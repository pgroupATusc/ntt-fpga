// NTT Accelerator

module NTT_Top #(
    parameter DATA_WIDTH_PER_INPUT = 28,
    parameter INPUT_PER_CYCLE = 64
  ) (
    inData,
    outData,
    in_start,
    out_start,
    clk,
    rst,
  );

  input clk, rst;

  input in_start[9:0];
  output logic out_start[9:0];

  input        [DATA_WIDTH_PER_INPUT-1:0] inData[INPUT_PER_CYCLE-1:0];
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_0_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_0_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_1_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_1_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_2_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_2_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_3_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_3_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_4_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_4_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_5_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_5_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_6_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_6_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_7_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_7_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_8_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_8_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_9_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_9_per_out[INPUT_PER_CYCLE-1:0];

  parameter [7:0] START_CYCLE[12] = {0, 7, 14, 21, 28, 35, 58, 82, 108, 138, 176, 230};

  // TODO(Tian): stage 0 32 butterfly units
  butterfly #(
    .start(START_CYCLE[0]),
    .factors({62736, 229351752, 248258143, 5986200, 141200910, 238271990, 210432655, 139336311,
              60410137, 227274721, 60657405, 217306794, 120438379, 125625707, 154088507, 162143577,
              168799557, 115574858, 163194978, 4369826, 90751938, 24738255, 174394830, 21511271,
              65612009, 151945076, 26268761, 224561048, 42684255, 135812431, 178512370, 96512966,
              8259075, 86907964, 229881708, 233570711, 81393489, 136863777, 184579826, 193086087,
              66137976, 46407972, 168246811, 9971642, 131575231, 215932086, 114248229, 132028761,
              104041706, 228870065, 39123511, 173212060, 110271140, 130565708, 151231163, 147718178,
              9497918, 131123953, 10785136, 167082925, 146990305, 12430538, 228578092, 263121861}))
  stage_0_butterfly_0 (
    .x_in(inData[0]),
    .y_in(inData[1]),
    .x_out(stage_0_per_in[0]),
    .y_out(stage_0_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({1907454, 18284087, 179300118, 3778321, 190023698, 215835949, 238852009, 79816727,
              90459251, 38780522, 188631715, 180949546, 93000404, 179673158, 68711843, 48588607,
              145932355, 25746466, 136072729, 68336365, 125408694, 31768873, 234613484, 42275209,
              18646649, 82056103, 241285957, 195819103, 249490832, 22776264, 138558999, 241947117,
              224650429, 132709741, 75771663, 106442355, 118813697, 213823426, 184231755, 222306946,
              48524018, 6841080, 184001594, 59811701, 149996455, 108455048, 9255299, 122257237,
              70352813, 244570986, 49444600, 48810421, 34248663, 35295690, 236243144, 231200794,
              125590824, 182424131, 135108737, 84704450, 176139969, 232516826, 129357001, 17124429}))
  stage_0_butterfly_1 (
    .x_in(inData[2]),
    .y_in(inData[3]),
    .x_out(stage_0_per_in[2]),
    .y_out(stage_0_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({127608977, 121332251, 157389868, 3052481, 238966374, 154495952, 172782070, 49806007,
              127870778, 70554670, 249304086, 54418504, 229943365, 135886727, 896607, 41484727,
              111929529, 235715975, 41726718, 27836602, 264371342, 149329993, 198700251, 228606302,
              140808004, 25249547, 155953488, 212109347, 105651651, 24888645, 95350060, 158561039,
              190509603, 260134415, 169809008, 236342274, 251686044, 130863524, 218474935, 244025737,
              65316150, 51724689, 179814135, 47156256, 122737973, 108348559, 239606434, 183216854,
              221042295, 267488469, 186854087, 198490305, 15301013, 97252224, 24230656, 109429555,
              104126955, 7378856, 72034061, 140793205, 83950689, 254596309, 184896958, 27247099}))
  stage_0_butterfly_2 (
    .x_in(inData[4]),
    .y_in(inData[5]),
    .x_out(stage_0_per_in[4]),
    .y_out(stage_0_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({169184935, 106831467, 195652857, 14448911, 91778054, 36311778, 32605484, 152480704,
              129584651, 110996066, 223960411, 45577523, 35630094, 68771072, 255719214, 48342959,
              123658638, 154830655, 202025824, 121686109, 210012123, 260828874, 140340588, 245765723,
              170942291, 125238212, 215941659, 20537000, 132315280, 129408474, 102742547, 44845193,
              180416915, 237936557, 30247571, 122360079, 104447750, 5132066, 197344625, 13810215,
              194219704, 162923321, 32737194, 103204044, 188122907, 217085295, 179717207, 92792804,
              72945707, 143112792, 210644544, 152283243, 249388588, 60682421, 181705475, 33223660,
              107928332, 119835732, 77051365, 150857390, 46671057, 122169973, 12667818, 34847782}))
  stage_0_butterfly_3 (
    .x_in(inData[6]),
    .y_in(inData[7]),
    .x_out(stage_0_per_in[6]),
    .y_out(stage_0_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({221849129, 151923798, 74962493, 133797910, 40496733, 2862602, 229751485, 117960054,
              173052617, 105948718, 254027033, 20059876, 200934478, 26464113, 77856633, 182951273,
              41023501, 34644106, 61497280, 265346073, 230823778, 131105010, 170978026, 44078325,
              132556999, 47307859, 24970434, 79305722, 136104512, 205576016, 61680409, 192247464,
              143100858, 233222120, 163860332, 134390440, 181610634, 153531059, 76430728, 101462472,
              181981633, 232770856, 98483239, 57501675, 207033531, 46461494, 228091235, 24794247,
              8255313, 238036964, 200339141, 59294895, 170921357, 118725672, 158126817, 110117913,
              38773847, 167554606, 171975768, 84361140, 247783732, 188917923, 69921988, 78030852}))
  stage_0_butterfly_4 (
    .x_in(inData[8]),
    .y_in(inData[9]),
    .x_out(stage_0_per_in[8]),
    .y_out(stage_0_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({172988180, 185050869, 67529023, 104771116, 41146808, 129899073, 88521257, 225676034,
              90342181, 243834156, 203523838, 156432226, 234989972, 116017893, 49058740, 247983171,
              51002920, 255155441, 18305869, 12986586, 67916891, 231410375, 225077819, 215954984,
              72252210, 112561771, 143573525, 227071465, 81013691, 119190794, 243451530, 60134449,
              124282928, 131237870, 198223, 249630983, 18803294, 201861189, 253464518, 107586283,
              129798040, 186098576, 185094855, 239753050, 265171130, 158309971, 160882583, 192193505,
              62374498, 219418748, 154596247, 32372991, 168351315, 33508832, 263412265, 106358666,
              118482368, 157437159, 248278309, 38642987, 26045295, 248241093, 36987199, 144111858}))
  stage_0_butterfly_5 (
    .x_in(inData[10]),
    .y_in(inData[11]),
    .x_out(stage_0_per_in[10]),
    .y_out(stage_0_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({163149532, 94277220, 144055138, 228780544, 120515996, 12984872, 55158081, 157537739,
              69936597, 63986967, 215111514, 171719097, 44459414, 184499901, 150205042, 152039665,
              227615757, 110912131, 246680455, 182209928, 6265971, 223045283, 110327668, 235787722,
              50475029, 36214289, 259992880, 14462331, 65760618, 54697818, 161245819, 259993096,
              87220148, 68196879, 39654333, 199075664, 81207363, 76114224, 7447708, 120912967,
              81762412, 106463701, 120134099, 227158983, 252263799, 170302338, 71887650, 228212013,
              122977291, 144673958, 519479, 123713876, 59384117, 178886927, 118024210, 199074208,
              110162160, 112635657, 79702710, 213908547, 17550542, 93347053, 132702632, 17823318}))
  stage_0_butterfly_6 (
    .x_in(inData[12]),
    .y_in(inData[13]),
    .x_out(stage_0_per_in[12]),
    .y_out(stage_0_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({196855462, 128643267, 205246482, 224318864, 131370540, 131972043, 68756958, 205821112,
              97670877, 34174616, 39872790, 265191298, 162528302, 51441041, 170882254, 171967455,
              138161289, 3764785, 200939178, 113870289, 234685655, 66804322, 210089549, 218637579,
              258291717, 92763586, 105582618, 222708254, 176214933, 234300746, 57174663, 259999423,
              7092568, 79425600, 37710032, 39822794, 267102876, 242814722, 145439741, 108148659,
              162088178, 194119116, 193601964, 28536923, 37647978, 57720967, 221029739, 195919352,
              7571096, 227038693, 23520122, 28811566, 225275209, 161625502, 164281505, 122116963,
              156290837, 185167965, 1058331, 117333915, 173307030, 193454786, 100165037, 83862241}))
  stage_0_butterfly_7 (
    .x_in(inData[14]),
    .y_in(inData[15]),
    .x_out(stage_0_per_in[14]),
    .y_out(stage_0_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({58836748, 155464901, 229152485, 255568559, 37016200, 757759, 30197592, 130707805,
              198671577, 137536510, 155288254, 237348335, 75750547, 141768337, 151080366, 223003866,
              24825033, 176371562, 244557461, 217608608, 164519211, 183965087, 98922830, 267382061,
              53079368, 49387461, 244197291, 64306041, 144216104, 30614038, 189539329, 119248989,
              215423485, 42144250, 99315902, 221060093, 196350608, 208391395, 206880652, 31181321,
              187622314, 169601951, 15282852, 131574531, 191761352, 68378584, 57198083, 146240700,
              228922625, 209673396, 245682235, 51270543, 149687609, 233335722, 135933105, 49462279,
              90978272, 8257788, 14827383, 212712674, 264868967, 239144038, 222406475, 126093548}))
  stage_0_butterfly_8 (
    .x_in(inData[16]),
    .y_in(inData[17]),
    .x_out(stage_0_per_in[16]),
    .y_out(stage_0_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({214715735, 235762007, 196177971, 205271224, 240473245, 211663060, 180175431, 109711544,
              238901161, 16804445, 199052238, 95429977, 56018142, 174653765, 99860276, 104275953,
              142361011, 214327170, 182231238, 39463122, 223844182, 260789685, 250127237, 130842873,
              231138525, 32828004, 247510253, 60661841, 150440065, 155312683, 158154241, 149391390,
              71354371, 230428614, 151814684, 106186088, 14667453, 69502239, 243146642, 215911494,
              58468223, 262471786, 94554508, 101824639, 250276575, 131432446, 215943874, 225035437,
              158081289, 192333550, 101905032, 8718982, 51995938, 15958207, 82860468, 71806036,
              264370556, 232696276, 235758123, 60363770, 103662145, 262883371, 183106668, 41823032}))
  stage_0_butterfly_9 (
    .x_in(inData[18]),
    .y_in(inData[19]),
    .x_out(stage_0_per_in[18]),
    .y_out(stage_0_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({102340758, 160425732, 129084525, 189138314, 183756330, 139937724, 57131388, 157541500,
              39614141, 225441652, 256641060, 97602587, 36695937, 190364932, 74424009, 43784819,
              173921335, 244546293, 233895150, 67840088, 237799186, 164954582, 252406953, 238836046,
              21531862, 62948694, 40943954, 110250618, 20254495, 109921777, 21576501, 123166625,
              164861991, 67538787, 70654895, 152866160, 101813716, 194581013, 152512971, 206403026,
              42011142, 250005524, 166506519, 224168732, 251811489, 138660240, 25877458, 14626898,
              181180691, 135180292, 94423638, 164438829, 147769827, 38284008, 115791483, 195002054,
              242430855, 195655909, 164243806, 5958674, 124253615, 192960909, 157152581, 219422045}))
  stage_0_butterfly_10 (
    .x_in(inData[20]),
    .y_in(inData[21]),
    .x_out(stage_0_per_in[20]),
    .y_out(stage_0_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({143786732, 75642576, 149881682, 257328955, 107655283, 234828316, 81142751, 174801883,
              159482341, 112432362, 134571988, 114891230, 110693156, 122092755, 185341670, 59653503,
              15577361, 229528882, 180088236, 76662541, 183904649, 159491283, 195538071, 204649844,
              256986339, 87947919, 255534095, 6777444, 45130170, 48856734, 129933587, 15637687,
              88993292, 81695275, 30549918, 261699407, 39931217, 237626776, 88157673, 190689455,
              259337446, 16392555, 51111850, 163665671, 256691758, 218881712, 107087275, 72197923,
              231263484, 243770087, 264251329, 48869357, 103488513, 202431138, 172857441, 99585718,
              11569899, 170722015, 164573784, 63257907, 158386056, 152845826, 65110284, 214283023}))
  stage_0_butterfly_11 (
    .x_in(inData[22]),
    .y_in(inData[23]),
    .x_out(stage_0_per_in[22]),
    .y_out(stage_0_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({98227373, 26796856, 29023980, 166961287, 161075491, 162545174, 23882789, 26873848,
              22558678, 264550106, 122229583, 157511077, 74718485, 246646236, 104073065, 103787038,
              128356119, 29220817, 38864951, 118901157, 178784227, 13711872, 173580392, 156914260,
              207607705, 198369788, 119226838, 240151518, 155144532, 95898316, 208507211, 148505031,
              239045807, 172925747, 154170583, 97938637, 84715346, 34838492, 2673613, 122693765,
              214985679, 61883556, 113130535, 65736109, 22397447, 231672458, 201302943, 110197348,
              220005950, 32796042, 241396543, 207300441, 174624298, 240095534, 77968856, 89434836,
              68807490, 49704806, 209917670, 221163181, 217428510, 117652871, 193565392, 86822274}))
  stage_0_butterfly_12 (
    .x_in(inData[24]),
    .y_in(inData[25]),
    .x_out(stage_0_per_in[24]),
    .y_out(stage_0_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({150057464, 192174913, 23448732, 205181101, 101070463, 200114, 63098068, 187534499,
              209153008, 188446087, 144072998, 77858155, 247373572, 78932104, 210239547, 268045200,
              122550241, 54047719, 183262830, 86866558, 71749872, 245038497, 180231688, 2963416,
              134429657, 113738086, 42021864, 247726047, 12808954, 77729422, 128052742, 212184418,
              126302082, 108404040, 6014167, 160990548, 78210348, 192227833, 252922274, 162344188,
              182834104, 225219172, 201087126, 239353906, 31027015, 127805784, 42785182, 259103093,
              33967221, 263029881, 48087349, 169234006, 181325168, 23443169, 139454911, 77508945,
              212592244, 240905155, 170346650, 51005918, 108779799, 83563004, 89733363, 193603540}))
  stage_0_butterfly_13 (
    .x_in(inData[26]),
    .y_in(inData[27]),
    .x_out(stage_0_per_in[26]),
    .y_out(stage_0_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({39962754, 83421235, 256558777, 14751178, 229530055, 110070131, 76671502, 71449616,
              260875356, 160647513, 10696564, 217600940, 25642441, 260649789, 109410131, 175074447,
              53554883, 114016424, 103692636, 213474870, 116165973, 179512630, 51440403, 188754097,
              266139878, 51323950, 216328989, 247259809, 173030765, 65690883, 114527376, 222486214,
              184347612, 116203844, 32820960, 33884144, 176100532, 5695672, 165433235, 140975706,
              163077087, 135684892, 89278624, 101029591, 256453055, 106059530, 149191288, 23651884,
              197994960, 119415929, 138451058, 141473040, 138996529, 26132679, 151037716, 12259140,
              49876629, 145011041, 220416699, 148939130, 1235353, 135766208, 183088464, 212842425}))
  stage_0_butterfly_14 (
    .x_in(inData[28]),
    .y_in(inData[29]),
    .x_out(stage_0_per_in[28]),
    .y_out(stage_0_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({93261610, 141812320, 172289773, 197944250, 254832984, 27854761, 258988459, 5510115,
              108081889, 126711917, 255307412, 59249925, 240106988, 86311355, 231600531, 103407625,
              159792872, 266701659, 94389433, 212384234, 126904432, 55935675, 211721600, 52557249,
              53728083, 205947916, 91288416, 50951254, 78692480, 154254400, 122077322, 56197115,
              16344528, 81573675, 88484653, 117319528, 187760701, 95352696, 132336250, 21476942,
              203097121, 80678005, 158896498, 21249308, 185758640, 258599303, 215878737, 114109699,
              39817818, 44100750, 36500136, 23918814, 34527937, 258759731, 116889475, 95430596,
              138868638, 11447146, 196733737, 103235635, 251183310, 180375437, 167274958, 58071796}))
  stage_0_butterfly_15 (
    .x_in(inData[30]),
    .y_in(inData[31]),
    .x_out(stage_0_per_in[30]),
    .y_out(stage_0_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({138390585, 232397550, 237695631, 76613625, 260020495, 251656189, 47407140, 30182006,
              50557363, 225306517, 63634221, 173443464, 126074738, 115237475, 131255494, 75233812,
              209093018, 85762236, 214996992, 59403344, 159528330, 174916329, 39518152, 238064453,
              221285249, 16499278, 71341164, 81430431, 171732518, 202855239, 73723002, 2615849,
              69789389, 1371159, 114463563, 196480564, 219691960, 139897823, 262334367, 199105134,
              229237307, 49661599, 253577157, 33454619, 127322073, 360580, 126370638, 85118780,
              103557733, 215247918, 187113601, 172102431, 55682893, 234938972, 256536575, 13664359,
              123998976, 18799530, 258162508, 242453874, 228964332, 197777956, 108727234, 261712272}))
  stage_0_butterfly_16 (
    .x_in(inData[32]),
    .y_in(inData[33]),
    .x_out(stage_0_per_in[32]),
    .y_out(stage_0_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({18568532, 173978412, 142538555, 183539945, 73697328, 35857213, 53030863, 202544817,
              148940015, 152136534, 148753884, 107281991, 35553140, 220692949, 249640388, 135453164,
              196709411, 145101039, 252862876, 56280600, 194605816, 236121751, 241597278, 254006109,
              121142478, 267007570, 206826789, 41756449, 147507351, 87928571, 240078055, 13493318,
              229741385, 21489734, 196341244, 187504892, 217792655, 247808775, 120846747, 28244848,
              86285917, 208868555, 182145624, 79440456, 48555419, 16609890, 2353936, 59625292,
              160793918, 1618864, 110273227, 205236559, 126498799, 46583536, 136554164, 99167958,
              57499821, 74632878, 53524475, 167937680, 86892569, 167199557, 244434992, 142049175}))
  stage_0_butterfly_17 (
    .x_in(inData[34]),
    .y_in(inData[35]),
    .x_out(stage_0_per_in[34]),
    .y_out(stage_0_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({5473511, 266521776, 144769477, 21572447, 46912433, 56987360, 26866408, 94223513,
              213245383, 20426733, 85422012, 66819851, 150130406, 181022773, 169515998, 203722503,
              132349487, 75105065, 221059178, 2011982, 11959677, 129605716, 219029055, 7229020,
              9479322, 206462525, 27115908, 234710989, 36246851, 107677384, 212385093, 194562323,
              130771778, 49717914, 163019788, 66144131, 107104549, 173951180, 107135677, 246477773,
              44515532, 251263130, 263884483, 185730304, 162829016, 14692215, 251425486, 255690434,
              87325743, 112251860, 211366667, 158126231, 86460683, 153141493, 151221429, 229582731,
              11703135, 100946881, 106563970, 34699254, 177264548, 149344309, 225116841, 151842442}))
  stage_0_butterfly_18 (
    .x_in(inData[36]),
    .y_in(inData[37]),
    .x_out(stage_0_per_in[36]),
    .y_out(stage_0_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({125480909, 184791819, 5231854, 151524267, 81083779, 56333048, 265950738, 179139190,
              81873483, 186348595, 4986407, 8297893, 155163691, 109371065, 208653574, 213678319,
              112142792, 174632895, 96892627, 258549338, 55192006, 194603131, 60603436, 28116292,
              155517338, 66449840, 260087354, 255738903, 90006293, 188542273, 242826313, 78592957,
              100132307, 5068353, 210363951, 96374025, 164529221, 29805745, 202640881, 197497401,
              256480283, 231677557, 123317306, 230350716, 6725515, 69230198, 218852619, 4491002,
              135171113, 116647317, 9249520, 244555167, 128889378, 90584256, 242671835, 47508483,
              48777982, 179869441, 30822536, 175007080, 188656071, 43714082, 56125789, 136274746}))
  stage_0_butterfly_19 (
    .x_in(inData[38]),
    .y_in(inData[39]),
    .x_out(stage_0_per_in[38]),
    .y_out(stage_0_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({234869713, 260851907, 226595737, 42776728, 206537906, 39521553, 189986560, 194846985,
              42053510, 15379209, 211444110, 61891902, 208159538, 254332699, 242184182, 192707093,
              234287689, 105706660, 76639397, 152738846, 228971558, 37752789, 245369685, 142898101,
              41652472, 158858535, 95816060, 145592959, 82875459, 185232992, 259733399, 204313060,
              186545936, 260923957, 261016176, 134614101, 243862110, 176789033, 112718220, 97251575,
              50106798, 13704349, 84901432, 222748125, 229222177, 109746000, 90105969, 263215622,
              266284483, 69414413, 148796874, 42275800, 135646873, 207530553, 148098547, 69218942,
              166068773, 53167918, 244602309, 150154963, 99177320, 110104975, 255918779, 57302073}))
  stage_0_butterfly_20 (
    .x_in(inData[40]),
    .y_in(inData[41]),
    .x_out(stage_0_per_in[40]),
    .y_out(stage_0_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({250606181, 29470818, 149138685, 54233307, 240784947, 132129988, 158533760, 248896168,
              212167090, 27029386, 228871862, 26659480, 205287356, 176832880, 61691447, 258883039,
              109505067, 21131779, 35559942, 66715025, 240649845, 229784592, 62782868, 115679885,
              159471860, 153682120, 235388028, 59375296, 230143339, 186483628, 143816111, 72475326,
              12651571, 157068444, 244905743, 54358169, 175334429, 260001724, 59370938, 209246609,
              58677377, 113781795, 249212399, 77840672, 225914175, 179365619, 38752877, 7116217,
              236327891, 263718984, 157430256, 158711864, 233906629, 74385386, 20877990, 198306293,
              220394580, 152365066, 198378776, 245615084, 265616179, 192872385, 260374016, 72549374}))
  stage_0_butterfly_21 (
    .x_in(inData[42]),
    .y_in(inData[43]),
    .x_out(stage_0_per_in[42]),
    .y_out(stage_0_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({5740730, 167586303, 218879515, 112058009, 116970950, 63216411, 104949331, 132200486,
              42733910, 83981669, 197423642, 12855237, 128505750, 171842488, 96976591, 96526884,
              151704879, 27233477, 154775650, 264329231, 109376139, 82632268, 162925843, 21764948,
              31551002, 144184457, 13842453, 235284227, 181725973, 83931467, 132907662, 97581367,
              63656435, 136382259, 230967163, 2029098, 149477651, 254244111, 185120393, 102116116,
              234954565, 227944808, 46729148, 89270439, 24734017, 213642756, 108647642, 212003953,
              150283834, 61250374, 67046513, 2557700, 136400329, 170944566, 28935497, 202918045,
              99410963, 206482017, 134843781, 235546264, 108704486, 117771098, 41112252, 220194496}))
  stage_0_butterfly_22 (
    .x_in(inData[44]),
    .y_in(inData[45]),
    .x_out(stage_0_per_in[44]),
    .y_out(stage_0_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({179625763, 148827249, 21458183, 1696019, 88419162, 58280814, 81930, 131559431,
              70436067, 192680584, 184608754, 13429213, 39140268, 39919904, 211152508, 115525972,
              234322267, 213843114, 111908324, 17233293, 243297654, 262250139, 78892295, 173572777,
              246940389, 162490819, 192516565, 82054424, 194815301, 108661782, 147106083, 157468594,
              88702124, 97492082, 59212137, 234121810, 159725962, 156378126, 145355888, 185671812,
              35430665, 164207528, 27694231, 78696193, 180249606, 204398753, 70151518, 99516991,
              21742303, 116801865, 212770879, 230635721, 106511467, 15750398, 171241703, 202001175,
              231268416, 130387641, 187415781, 37225330, 138920976, 18191490, 179287997, 159562860}))
  stage_0_butterfly_23 (
    .x_in(inData[46]),
    .y_in(inData[47]),
    .x_out(stage_0_per_in[46]),
    .y_out(stage_0_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({106056773, 48491280, 208950205, 6668530, 239404299, 24825329, 263982663, 185532067,
              240039943, 136783171, 57437223, 211688613, 100943177, 209177739, 4470762, 41306715,
              136599943, 24132582, 18792168, 146607869, 179831843, 111072250, 212470099, 208828758,
              7369182, 171197489, 144151142, 168472713, 116861206, 58714599, 134997518, 206941931,
              50402804, 183351284, 45294283, 44427932, 124269051, 233581580, 168938760, 130959181,
              159543175, 215737735, 25904197, 84557377, 223537938, 165004785, 151696189, 10658994,
              106146355, 7620297, 213752765, 223629100, 3104477, 165252821, 204917473, 38635824,
              152734723, 264133989, 89201641, 76772605, 10598408, 141503129, 164702238, 166754761}))
  stage_0_butterfly_24 (
    .x_in(inData[48]),
    .y_in(inData[49]),
    .x_out(stage_0_per_in[48]),
    .y_out(stage_0_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({58136368, 268021045, 201838233, 155885829, 170979076, 194935198, 63162591, 103408097,
              83840449, 216659963, 248573392, 190439637, 225546029, 155010430, 15349425, 239742054,
              177927774, 66663233, 201356021, 179809501, 113458040, 201979579, 6044206, 206641346,
              184067420, 127364429, 70489814, 14129846, 136415646, 53126633, 204076371, 134053105,
              118651137, 111920700, 98566622, 132259857, 125694138, 231794807, 107070533, 157805049,
              250060684, 227465231, 90061976, 27951846, 47826324, 168435324, 226717406, 246208472,
              61116726, 235669313, 120964758, 52189384, 136046821, 40354434, 165567634, 131200140,
              169435715, 203745198, 24603905, 13532798, 123887389, 237430063, 55517835, 23085612}))
  stage_0_butterfly_25 (
    .x_in(inData[50]),
    .y_in(inData[51]),
    .x_out(stage_0_per_in[50]),
    .y_out(stage_0_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({104423755, 68227492, 189611269, 73017801, 21594518, 9880764, 225369254, 156474406,
              264479828, 127467506, 16955107, 169350110, 183488163, 32128041, 179315380, 60805498,
              27503451, 52676293, 171672871, 83253386, 122367942, 172273878, 104310584, 223368694,
              33019077, 83749497, 156153949, 56381879, 241508336, 138905259, 205242093, 221722750,
              195906424, 107691461, 9245191, 51218933, 184151583, 137830340, 236547476, 232729335,
              67287217, 195074984, 129666909, 4952604, 172140914, 16462324, 176366269, 55752506,
              188909348, 253757449, 230339059, 73689066, 16063721, 169231043, 54766528, 205614247,
              241821884, 95072757, 254310437, 264371786, 210853880, 230124651, 221585216, 207505578}))
  stage_0_butterfly_26 (
    .x_in(inData[52]),
    .y_in(inData[53]),
    .x_out(stage_0_per_in[52]),
    .y_out(stage_0_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({136664320, 135770551, 224508026, 92074820, 92366490, 203810197, 78969227, 91588944,
              139852785, 62704870, 204252016, 236052416, 106354792, 259685293, 168672066, 171138130,
              81860583, 134876482, 111274912, 55730854, 133008104, 152468473, 99112512, 26767263,
              99821278, 92092447, 34336755, 168849030, 216240230, 87141435, 69177824, 96021565,
              181033780, 201880574, 59669292, 160584715, 245310720, 2176252, 138198441, 248617642,
              106129670, 180394230, 101060936, 229121016, 105408561, 171482266, 129184142, 183002860,
              194876189, 40301047, 74816213, 73137377, 71660202, 28921814, 185723977, 152308098,
              205958875, 30940476, 83294274, 154688443, 242290819, 144681042, 163860385, 234273255}))
  stage_0_butterfly_27 (
    .x_in(inData[54]),
    .y_in(inData[55]),
    .x_out(stage_0_per_in[54]),
    .y_out(stage_0_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({63355713, 198563101, 224551623, 244373783, 89303497, 198839540, 59001681, 227953669,
              265709143, 135413478, 58605619, 118174461, 6291440, 36389566, 146899744, 213475348,
              260400385, 245230909, 209546662, 170534402, 184276602, 158032303, 234070704, 190758660,
              102903513, 115048608, 224670583, 203514552, 45907501, 62285640, 56939589, 150485586,
              65941195, 43314683, 93988508, 265006255, 68363059, 197478524, 19830371, 110482921,
              85558096, 67824335, 141580746, 135142897, 98503463, 174146267, 160170338, 183449518,
              79129285, 96257044, 124727876, 218509565, 291007, 227652594, 255492938, 148811231,
              237882452, 74916156, 8009648, 251093184, 127215407, 140577689, 83000954, 34079608}))
  stage_0_butterfly_28 (
    .x_in(inData[56]),
    .y_in(inData[57]),
    .x_out(stage_0_per_in[56]),
    .y_out(stage_0_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({101375441, 95052731, 83959851, 112531453, 142276463, 85927424, 228944741, 215784466,
              147276523, 167238213, 175168807, 230885966, 22914950, 196216182, 137992276, 19847969,
              130985550, 249112263, 198284911, 215285662, 175012394, 178662179, 152315952, 154802450,
              118213444, 40802701, 4622329, 201888697, 153503748, 113731328, 225486456, 68532350,
              107657151, 200590842, 216371534, 255059903, 136530068, 214972665, 35417568, 202258967,
              105733032, 23130727, 7430278, 246714101, 41771488, 208345113, 30147565, 23277706,
              258487225, 117177606, 32948426, 57795922, 177554441, 161226237, 68094050, 82689315,
              149425076, 195813478, 117454680, 44226281, 82939526, 208881897, 117458270, 171515704}))
  stage_0_butterfly_29 (
    .x_in(inData[58]),
    .y_in(inData[59]),
    .x_out(stage_0_per_in[58]),
    .y_out(stage_0_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({173776705, 37560959, 130521421, 218305863, 149796825, 37761143, 167654012, 25592978,
              69963660, 177400482, 242086614, 125945553, 154162735, 88343680, 163943008, 41373747,
              96784305, 27425418, 178609958, 99694466, 183166375, 239054686, 264712232, 137079211,
              42583023, 177007616, 237453043, 237567768, 68847542, 200029177, 245228415, 257632808,
              17252496, 236356015, 20606850, 148722321, 97520605, 50703780, 151289170, 113484891,
              111517965, 26760307, 41328094, 11562888, 140190159, 224658359, 82596723, 130055322,
              268107376, 625780, 92713113, 215495577, 217198560, 89497967, 44239577, 211488291,
              163847221, 216947907, 13484173, 246176063, 48025256, 42743336, 95081716, 76694868}))
  stage_0_butterfly_30 (
    .x_in(inData[60]),
    .y_in(inData[61]),
    .x_out(stage_0_per_in[60]),
    .y_out(stage_0_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({99627052, 17746678, 36284828, 145182880, 193094875, 235736575, 106508361, 228413454,
              178085825, 10710243, 67348921, 216347827, 120761900, 45256937, 247160596, 32751373,
              150225643, 143680187, 241625831, 192995301, 139998882, 168382927, 267141235, 139421138,
              249903585, 209077448, 259081121, 103000049, 134859556, 3595020, 163361339, 99532395,
              26620819, 134045502, 32461064, 83014713, 98179318, 91252917, 213289884, 250977019,
              226850270, 17172477, 68554215, 101673356, 216246538, 161740894, 124135460, 90052819,
              74278900, 17691838, 97283065, 266251087, 118163582, 213947035, 159360601, 134709760,
              192889387, 1741916, 65815578, 45566469, 58580381, 107220558, 239548624, 127926589}))
  stage_0_butterfly_31 (
    .x_in(inData[62]),
    .y_in(inData[63]),
    .x_out(stage_0_per_in[62]),
    .y_out(stage_0_per_in[63]),
    .clk(clk),
    .rst(rst)
  );





  // TODO(Yang): stage 0 -> stage 1 permutation
  // FIXME: ignore butterfly units for now.
  stage_0_permutation #(
    .DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    .INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_0_1_per (
    .inData_0(stage_0_per_in[0]),
    .inData_1(stage_0_per_in[1]),
    .inData_2(stage_0_per_in[2]),
    .inData_3(stage_0_per_in[3]),
    .inData_4(stage_0_per_in[4]),
    .inData_5(stage_0_per_in[5]),
    .inData_6(stage_0_per_in[6]),
    .inData_7(stage_0_per_in[7]),
    .inData_8(stage_0_per_in[8]),
    .inData_9(stage_0_per_in[9]),
    .inData_10(stage_0_per_in[10]),
    .inData_11(stage_0_per_in[11]),
    .inData_12(stage_0_per_in[12]),
    .inData_13(stage_0_per_in[13]),
    .inData_14(stage_0_per_in[14]),
    .inData_15(stage_0_per_in[15]),
    .inData_16(stage_0_per_in[16]),
    .inData_17(stage_0_per_in[17]),
    .inData_18(stage_0_per_in[18]),
    .inData_19(stage_0_per_in[19]),
    .inData_20(stage_0_per_in[20]),
    .inData_21(stage_0_per_in[21]),
    .inData_22(stage_0_per_in[22]),
    .inData_23(stage_0_per_in[23]),
    .inData_24(stage_0_per_in[24]),
    .inData_25(stage_0_per_in[25]),
    .inData_26(stage_0_per_in[26]),
    .inData_27(stage_0_per_in[27]),
    .inData_28(stage_0_per_in[28]),
    .inData_29(stage_0_per_in[29]),
    .inData_30(stage_0_per_in[30]),
    .inData_31(stage_0_per_in[31]),
    .inData_32(stage_0_per_in[32]),
    .inData_33(stage_0_per_in[33]),
    .inData_34(stage_0_per_in[34]),
    .inData_35(stage_0_per_in[35]),
    .inData_36(stage_0_per_in[36]),
    .inData_37(stage_0_per_in[37]),
    .inData_38(stage_0_per_in[38]),
    .inData_39(stage_0_per_in[39]),
    .inData_40(stage_0_per_in[40]),
    .inData_41(stage_0_per_in[41]),
    .inData_42(stage_0_per_in[42]),
    .inData_43(stage_0_per_in[43]),
    .inData_44(stage_0_per_in[44]),
    .inData_45(stage_0_per_in[45]),
    .inData_46(stage_0_per_in[46]),
    .inData_47(stage_0_per_in[47]),
    .inData_48(stage_0_per_in[48]),
    .inData_49(stage_0_per_in[49]),
    .inData_50(stage_0_per_in[50]),
    .inData_51(stage_0_per_in[51]),
    .inData_52(stage_0_per_in[52]),
    .inData_53(stage_0_per_in[53]),
    .inData_54(stage_0_per_in[54]),
    .inData_55(stage_0_per_in[55]),
    .inData_56(stage_0_per_in[56]),
    .inData_57(stage_0_per_in[57]),
    .inData_58(stage_0_per_in[58]),
    .inData_59(stage_0_per_in[59]),
    .inData_60(stage_0_per_in[60]),
    .inData_61(stage_0_per_in[61]),
    .inData_62(stage_0_per_in[62]),
    .inData_63(stage_0_per_in[63]),
    .outData_0(stage_0_per_out[0]),
    .outData_1(stage_0_per_out[1]),
    .outData_2(stage_0_per_out[2]),
    .outData_3(stage_0_per_out[3]),
    .outData_4(stage_0_per_out[4]),
    .outData_5(stage_0_per_out[5]),
    .outData_6(stage_0_per_out[6]),
    .outData_7(stage_0_per_out[7]),
    .outData_8(stage_0_per_out[8]),
    .outData_9(stage_0_per_out[9]),
    .outData_10(stage_0_per_out[10]),
    .outData_11(stage_0_per_out[11]),
    .outData_12(stage_0_per_out[12]),
    .outData_13(stage_0_per_out[13]),
    .outData_14(stage_0_per_out[14]),
    .outData_15(stage_0_per_out[15]),
    .outData_16(stage_0_per_out[16]),
    .outData_17(stage_0_per_out[17]),
    .outData_18(stage_0_per_out[18]),
    .outData_19(stage_0_per_out[19]),
    .outData_20(stage_0_per_out[20]),
    .outData_21(stage_0_per_out[21]),
    .outData_22(stage_0_per_out[22]),
    .outData_23(stage_0_per_out[23]),
    .outData_24(stage_0_per_out[24]),
    .outData_25(stage_0_per_out[25]),
    .outData_26(stage_0_per_out[26]),
    .outData_27(stage_0_per_out[27]),
    .outData_28(stage_0_per_out[28]),
    .outData_29(stage_0_per_out[29]),
    .outData_30(stage_0_per_out[30]),
    .outData_31(stage_0_per_out[31]),
    .outData_32(stage_0_per_out[32]),
    .outData_33(stage_0_per_out[33]),
    .outData_34(stage_0_per_out[34]),
    .outData_35(stage_0_per_out[35]),
    .outData_36(stage_0_per_out[36]),
    .outData_37(stage_0_per_out[37]),
    .outData_38(stage_0_per_out[38]),
    .outData_39(stage_0_per_out[39]),
    .outData_40(stage_0_per_out[40]),
    .outData_41(stage_0_per_out[41]),
    .outData_42(stage_0_per_out[42]),
    .outData_43(stage_0_per_out[43]),
    .outData_44(stage_0_per_out[44]),
    .outData_45(stage_0_per_out[45]),
    .outData_46(stage_0_per_out[46]),
    .outData_47(stage_0_per_out[47]),
    .outData_48(stage_0_per_out[48]),
    .outData_49(stage_0_per_out[49]),
    .outData_50(stage_0_per_out[50]),
    .outData_51(stage_0_per_out[51]),
    .outData_52(stage_0_per_out[52]),
    .outData_53(stage_0_per_out[53]),
    .outData_54(stage_0_per_out[54]),
    .outData_55(stage_0_per_out[55]),
    .outData_56(stage_0_per_out[56]),
    .outData_57(stage_0_per_out[57]),
    .outData_58(stage_0_per_out[58]),
    .outData_59(stage_0_per_out[59]),
    .outData_60(stage_0_per_out[60]),
    .outData_61(stage_0_per_out[61]),
    .outData_62(stage_0_per_out[62]),
    .outData_63(stage_0_per_out[63]),
    .in_start(in_start[0]),
    .out_start(out_start[0]),
    .clk(clk),
    .rst(rst)
  );

  // TODO(Tian): stage 1 32 butterfly units
  butterfly #(
    .start(START_CYCLE[1]),
    .factors({178626802, 36426289, 226568978, 228368554, 142863934, 98446051, 100723721, 195462811,
              25937392, 48496256, 26964940, 236960516, 49890248, 58870518, 57740084, 148535761,
              238700391, 170998790, 81363847, 54281363, 185850221, 153913781, 35411505, 90710559,
              135389110, 26451456, 34884345, 189299702, 212020732, 50385541, 214331009, 46629005,
              200295213, 6208689, 154135831, 99461488, 156023579, 47430573, 139714595, 143466178,
              214078274, 118216948, 264282458, 173116375, 197485473, 9453674, 167134668, 157049837,
              245518247, 43737855, 195063937, 264289232, 205675156, 54092187, 251274354, 198072981,
              44349942, 100770703, 120419308, 224620084, 75240990, 267404879, 143647295, 133881133}))
  stage_1_butterfly_0 (
    .x_in(stage_0_per_out[0]),
    .y_in(stage_0_per_out[1]),
    .x_out(stage_1_per_in[0]),
    .y_out(stage_1_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({178626802, 36426289, 226568978, 228368554, 142863934, 98446051, 100723721, 195462811,
              25937392, 48496256, 26964940, 236960516, 49890248, 58870518, 57740084, 148535761,
              238700391, 170998790, 81363847, 54281363, 185850221, 153913781, 35411505, 90710559,
              135389110, 26451456, 34884345, 189299702, 212020732, 50385541, 214331009, 46629005,
              200295213, 6208689, 154135831, 99461488, 156023579, 47430573, 139714595, 143466178,
              214078274, 118216948, 264282458, 173116375, 197485473, 9453674, 167134668, 157049837,
              245518247, 43737855, 195063937, 264289232, 205675156, 54092187, 251274354, 198072981,
              44349942, 100770703, 120419308, 224620084, 75240990, 267404879, 143647295, 133881133}))
  stage_1_butterfly_1 (
    .x_in(stage_0_per_out[2]),
    .y_in(stage_0_per_out[3]),
    .x_out(stage_1_per_in[2]),
    .y_out(stage_1_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({241419299, 189966412, 57439678, 104968162, 115334054, 213018760, 66106013, 150529015,
              66456987, 266940341, 79732409, 61436946, 185097589, 230680452, 136199054, 72619804,
              101221270, 65241583, 161494327, 129726580, 227605745, 196403691, 3059556, 262108538,
              111262804, 39377609, 170188367, 188624074, 148511346, 175901771, 109286034, 124518160,
              40738286, 39161232, 180106398, 219432305, 79909455, 259358426, 209076586, 145040924,
              107222748, 106026444, 136983182, 119641299, 231584900, 118804291, 145952502, 58085086,
              260055946, 26707009, 268223107, 141552463, 178774268, 68124275, 5742112, 73785583,
              186303790, 89556414, 90238900, 211474022, 135620074, 80152118, 59970273, 78067214}))
  stage_1_butterfly_2 (
    .x_in(stage_0_per_out[4]),
    .y_in(stage_0_per_out[5]),
    .x_out(stage_1_per_in[4]),
    .y_out(stage_1_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({241419299, 189966412, 57439678, 104968162, 115334054, 213018760, 66106013, 150529015,
              66456987, 266940341, 79732409, 61436946, 185097589, 230680452, 136199054, 72619804,
              101221270, 65241583, 161494327, 129726580, 227605745, 196403691, 3059556, 262108538,
              111262804, 39377609, 170188367, 188624074, 148511346, 175901771, 109286034, 124518160,
              40738286, 39161232, 180106398, 219432305, 79909455, 259358426, 209076586, 145040924,
              107222748, 106026444, 136983182, 119641299, 231584900, 118804291, 145952502, 58085086,
              260055946, 26707009, 268223107, 141552463, 178774268, 68124275, 5742112, 73785583,
              186303790, 89556414, 90238900, 211474022, 135620074, 80152118, 59970273, 78067214}))
  stage_1_butterfly_3 (
    .x_in(stage_0_per_out[6]),
    .y_in(stage_0_per_out[7]),
    .x_out(stage_1_per_in[6]),
    .y_out(stage_1_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({202037642, 141057137, 124029413, 258951073, 144625416, 83042590, 152694343, 247893310,
              113912362, 153843002, 9977836, 203299319, 194834330, 127868408, 267034870, 90431622,
              255819997, 190155959, 92670067, 25148713, 10513337, 224762304, 65501903, 72006316,
              38583127, 138773321, 219164507, 34739971, 160223263, 60791061, 202709135, 154200425,
              111948379, 248800534, 158020658, 20654843, 87171014, 84553412, 73987125, 89839882,
              71023991, 208367077, 109238580, 140702439, 144486207, 198469359, 156384032, 243002151,
              66619308, 255369977, 136306850, 27101256, 204183192, 215044990, 37830528, 176150397,
              230038199, 84103703, 37832342, 109081133, 184194991, 161356640, 85850918, 61148806}))
  stage_1_butterfly_4 (
    .x_in(stage_0_per_out[8]),
    .y_in(stage_0_per_out[9]),
    .x_out(stage_1_per_in[8]),
    .y_out(stage_1_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({202037642, 141057137, 124029413, 258951073, 144625416, 83042590, 152694343, 247893310,
              113912362, 153843002, 9977836, 203299319, 194834330, 127868408, 267034870, 90431622,
              255819997, 190155959, 92670067, 25148713, 10513337, 224762304, 65501903, 72006316,
              38583127, 138773321, 219164507, 34739971, 160223263, 60791061, 202709135, 154200425,
              111948379, 248800534, 158020658, 20654843, 87171014, 84553412, 73987125, 89839882,
              71023991, 208367077, 109238580, 140702439, 144486207, 198469359, 156384032, 243002151,
              66619308, 255369977, 136306850, 27101256, 204183192, 215044990, 37830528, 176150397,
              230038199, 84103703, 37832342, 109081133, 184194991, 161356640, 85850918, 61148806}))
  stage_1_butterfly_5 (
    .x_in(stage_0_per_out[10]),
    .y_in(stage_0_per_out[11]),
    .x_out(stage_1_per_in[10]),
    .y_out(stage_1_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({224076531, 75414331, 176876579, 55709426, 42559975, 9179161, 181657279, 95442771,
              179710610, 188476710, 131815160, 214979600, 22106362, 127510598, 251982020, 217412044,
              161018204, 82911469, 54856389, 34957318, 141500462, 176271587, 138344594, 207338429,
              36505175, 35544064, 107122996, 89363633, 183471966, 79351768, 263768524, 245466834,
              79007221, 72719897, 75051406, 104015737, 254205318, 77136822, 48961458, 73243528,
              236016875, 16967674, 41046131, 205950205, 263500442, 20490089, 238066757, 176574100,
              173525016, 215608734, 146660836, 207179347, 2306944, 217413665, 233611200, 76831465,
              249749550, 131659808, 111544693, 252140774, 216035935, 201376724, 86146205, 115561740}))
  stage_1_butterfly_6 (
    .x_in(stage_0_per_out[12]),
    .y_in(stage_0_per_out[13]),
    .x_out(stage_1_per_in[12]),
    .y_out(stage_1_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({224076531, 75414331, 176876579, 55709426, 42559975, 9179161, 181657279, 95442771,
              179710610, 188476710, 131815160, 214979600, 22106362, 127510598, 251982020, 217412044,
              161018204, 82911469, 54856389, 34957318, 141500462, 176271587, 138344594, 207338429,
              36505175, 35544064, 107122996, 89363633, 183471966, 79351768, 263768524, 245466834,
              79007221, 72719897, 75051406, 104015737, 254205318, 77136822, 48961458, 73243528,
              236016875, 16967674, 41046131, 205950205, 263500442, 20490089, 238066757, 176574100,
              173525016, 215608734, 146660836, 207179347, 2306944, 217413665, 233611200, 76831465,
              249749550, 131659808, 111544693, 252140774, 216035935, 201376724, 86146205, 115561740}))
  stage_1_butterfly_7 (
    .x_in(stage_0_per_out[14]),
    .y_in(stage_0_per_out[15]),
    .x_out(stage_1_per_in[14]),
    .y_out(stage_1_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({262853884, 204172184, 202016934, 144194814, 200835165, 155441062, 139662643, 209967729,
              213369302, 193915015, 48721923, 222818810, 77445892, 151896708, 41376169, 207289252,
              260565899, 192679930, 80939041, 40189829, 28923545, 169229772, 89821167, 74346844,
              221852517, 216420108, 116261862, 150921330, 81165688, 172134458, 254651521, 143985240,
              251186267, 188623776, 173013758, 192273850, 7373784, 202075477, 33406019, 76213351,
              256339290, 259641163, 2568552, 94417879, 66687, 82259521, 14131216, 226423252,
              117147237, 259932536, 2885885, 232035425, 69918547, 166849602, 13809973, 217984510,
              195258296, 144316291, 232016200, 91036891, 224618046, 18026307, 24281843, 168335279}))
  stage_1_butterfly_8 (
    .x_in(stage_0_per_out[16]),
    .y_in(stage_0_per_out[17]),
    .x_out(stage_1_per_in[16]),
    .y_out(stage_1_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({262853884, 204172184, 202016934, 144194814, 200835165, 155441062, 139662643, 209967729,
              213369302, 193915015, 48721923, 222818810, 77445892, 151896708, 41376169, 207289252,
              260565899, 192679930, 80939041, 40189829, 28923545, 169229772, 89821167, 74346844,
              221852517, 216420108, 116261862, 150921330, 81165688, 172134458, 254651521, 143985240,
              251186267, 188623776, 173013758, 192273850, 7373784, 202075477, 33406019, 76213351,
              256339290, 259641163, 2568552, 94417879, 66687, 82259521, 14131216, 226423252,
              117147237, 259932536, 2885885, 232035425, 69918547, 166849602, 13809973, 217984510,
              195258296, 144316291, 232016200, 91036891, 224618046, 18026307, 24281843, 168335279}))
  stage_1_butterfly_9 (
    .x_in(stage_0_per_out[18]),
    .y_in(stage_0_per_out[19]),
    .x_out(stage_1_per_in[18]),
    .y_out(stage_1_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({243595082, 114289273, 205274966, 80852279, 13214022, 183986337, 4628244, 255259435,
              204246510, 146691665, 27222642, 165177241, 90803899, 253065021, 156486669, 182882105,
              2705617, 171586403, 94113816, 154399218, 35769351, 177621090, 180859208, 27789608,
              234383020, 103427147, 37907807, 180135303, 82858612, 111988251, 67895486, 75455626,
              212990958, 176645554, 239438610, 244247525, 82105625, 197737960, 223749061, 204890405,
              193207980, 258770065, 22039584, 7487276, 198659369, 149046252, 33154381, 33861678,
              46680870, 64324001, 57534183, 212068395, 197375798, 248421583, 211651639, 262436297,
              85354678, 239135625, 230913482, 186920055, 242981970, 119165597, 118812967, 88850354}))
  stage_1_butterfly_10 (
    .x_in(stage_0_per_out[20]),
    .y_in(stage_0_per_out[21]),
    .x_out(stage_1_per_in[20]),
    .y_out(stage_1_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({243595082, 114289273, 205274966, 80852279, 13214022, 183986337, 4628244, 255259435,
              204246510, 146691665, 27222642, 165177241, 90803899, 253065021, 156486669, 182882105,
              2705617, 171586403, 94113816, 154399218, 35769351, 177621090, 180859208, 27789608,
              234383020, 103427147, 37907807, 180135303, 82858612, 111988251, 67895486, 75455626,
              212990958, 176645554, 239438610, 244247525, 82105625, 197737960, 223749061, 204890405,
              193207980, 258770065, 22039584, 7487276, 198659369, 149046252, 33154381, 33861678,
              46680870, 64324001, 57534183, 212068395, 197375798, 248421583, 211651639, 262436297,
              85354678, 239135625, 230913482, 186920055, 242981970, 119165597, 118812967, 88850354}))
  stage_1_butterfly_11 (
    .x_in(stage_0_per_out[22]),
    .y_in(stage_0_per_out[23]),
    .x_out(stage_1_per_in[22]),
    .y_out(stage_1_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({256992454, 266373219, 239354922, 34279912, 86047893, 209875154, 84463383, 121172029,
              174110644, 250769297, 116219557, 242437879, 35608242, 181957723, 28513237, 25651112,
              230880884, 207436891, 9083394, 35697312, 254464819, 29380441, 63900610, 34535827,
              37207751, 104305160, 259466327, 22230677, 258848760, 245673827, 225061179, 211697180,
              7004663, 154780521, 156508649, 76495986, 193530415, 113066699, 173627934, 112847505,
              208392312, 139316176, 161193348, 184571212, 256317058, 178875242, 96851793, 247989601,
              104721465, 155494097, 188253439, 147907047, 194631063, 243436973, 218464636, 177240151,
              175705236, 138028127, 144500142, 106663692, 250268531, 110007683, 208182039, 78372181}))
  stage_1_butterfly_12 (
    .x_in(stage_0_per_out[24]),
    .y_in(stage_0_per_out[25]),
    .x_out(stage_1_per_in[24]),
    .y_out(stage_1_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({256992454, 266373219, 239354922, 34279912, 86047893, 209875154, 84463383, 121172029,
              174110644, 250769297, 116219557, 242437879, 35608242, 181957723, 28513237, 25651112,
              230880884, 207436891, 9083394, 35697312, 254464819, 29380441, 63900610, 34535827,
              37207751, 104305160, 259466327, 22230677, 258848760, 245673827, 225061179, 211697180,
              7004663, 154780521, 156508649, 76495986, 193530415, 113066699, 173627934, 112847505,
              208392312, 139316176, 161193348, 184571212, 256317058, 178875242, 96851793, 247989601,
              104721465, 155494097, 188253439, 147907047, 194631063, 243436973, 218464636, 177240151,
              175705236, 138028127, 144500142, 106663692, 250268531, 110007683, 208182039, 78372181}))
  stage_1_butterfly_13 (
    .x_in(stage_0_per_out[26]),
    .y_in(stage_0_per_out[27]),
    .x_out(stage_1_per_in[26]),
    .y_out(stage_1_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({77239454, 148884778, 143734200, 236741674, 222855093, 57044952, 86334506, 126959268,
              21923530, 126650083, 186026798, 33343400, 26776855, 40931981, 42903438, 63912782,
              58103200, 166350047, 239780428, 91136142, 251689720, 110850189, 253128696, 81924749,
              197145719, 187446019, 56848151, 255364493, 164222678, 124441328, 79432680, 39292866,
              143288167, 210949816, 22021280, 117619035, 248341796, 123481104, 27523605, 153827860,
              197016099, 250734390, 171258656, 106713399, 262755833, 108936038, 60493834, 152193297,
              13327732, 130184658, 14594411, 260941520, 193102647, 267667077, 218565763, 162889363,
              57880935, 98151275, 202657965, 141192231, 145663803, 142379740, 68372869, 252921174}))
  stage_1_butterfly_14 (
    .x_in(stage_0_per_out[28]),
    .y_in(stage_0_per_out[29]),
    .x_out(stage_1_per_in[28]),
    .y_out(stage_1_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({77239454, 148884778, 143734200, 236741674, 222855093, 57044952, 86334506, 126959268,
              21923530, 126650083, 186026798, 33343400, 26776855, 40931981, 42903438, 63912782,
              58103200, 166350047, 239780428, 91136142, 251689720, 110850189, 253128696, 81924749,
              197145719, 187446019, 56848151, 255364493, 164222678, 124441328, 79432680, 39292866,
              143288167, 210949816, 22021280, 117619035, 248341796, 123481104, 27523605, 153827860,
              197016099, 250734390, 171258656, 106713399, 262755833, 108936038, 60493834, 152193297,
              13327732, 130184658, 14594411, 260941520, 193102647, 267667077, 218565763, 162889363,
              57880935, 98151275, 202657965, 141192231, 145663803, 142379740, 68372869, 252921174}))
  stage_1_butterfly_15 (
    .x_in(stage_0_per_out[30]),
    .y_in(stage_0_per_out[31]),
    .x_out(stage_1_per_in[30]),
    .y_out(stage_1_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({22329094, 150629496, 146360154, 175887545, 70370832, 171269635, 124927121, 236561162,
              43396787, 213843220, 37292607, 91188581, 52859373, 108521058, 41918325, 67911621,
              224183590, 104486975, 129161289, 100791881, 67400723, 247062782, 48447796, 211284483,
              260125445, 46126435, 199208092, 222236846, 157341419, 31157387, 246555646, 38115064,
              72618725, 145706676, 222840723, 106939991, 116859647, 264758616, 184120139, 17337072,
              38429557, 195763450, 253615348, 3677235, 236609676, 126894636, 19066791, 66528431,
              53251080, 179997990, 41015351, 81431484, 64307891, 204816575, 167135704, 91524025,
              254723792, 75117738, 147133292, 141917139, 4884476, 254692251, 124656108, 45684920}))
  stage_1_butterfly_16 (
    .x_in(stage_0_per_out[32]),
    .y_in(stage_0_per_out[33]),
    .x_out(stage_1_per_in[32]),
    .y_out(stage_1_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({22329094, 150629496, 146360154, 175887545, 70370832, 171269635, 124927121, 236561162,
              43396787, 213843220, 37292607, 91188581, 52859373, 108521058, 41918325, 67911621,
              224183590, 104486975, 129161289, 100791881, 67400723, 247062782, 48447796, 211284483,
              260125445, 46126435, 199208092, 222236846, 157341419, 31157387, 246555646, 38115064,
              72618725, 145706676, 222840723, 106939991, 116859647, 264758616, 184120139, 17337072,
              38429557, 195763450, 253615348, 3677235, 236609676, 126894636, 19066791, 66528431,
              53251080, 179997990, 41015351, 81431484, 64307891, 204816575, 167135704, 91524025,
              254723792, 75117738, 147133292, 141917139, 4884476, 254692251, 124656108, 45684920}))
  stage_1_butterfly_17 (
    .x_in(stage_0_per_out[34]),
    .y_in(stage_0_per_out[35]),
    .x_out(stage_1_per_in[34]),
    .y_out(stage_1_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({114906207, 95956458, 93815079, 119248786, 244981517, 25402945, 164849679, 253446904,
              182759226, 65939487, 218411001, 105651679, 13136617, 86425411, 248430418, 104273059,
              48258409, 32326785, 86611832, 248049881, 220409117, 60951044, 98839404, 128923754,
              50041017, 51590619, 71466452, 81879124, 6839312, 50250252, 70993112, 202017141,
              77785137, 166705511, 159555178, 176106545, 168682489, 99151986, 45900567, 135965343,
              95745785, 196552678, 266184237, 36678208, 124689641, 250979164, 196076822, 242448751,
              142932928, 232700332, 26885190, 157159811, 187973069, 49412866, 195777196, 24169593,
              242906033, 123556687, 258128862, 66398989, 60114085, 79759830, 203861878, 47380903}))
  stage_1_butterfly_18 (
    .x_in(stage_0_per_out[36]),
    .y_in(stage_0_per_out[37]),
    .x_out(stage_1_per_in[36]),
    .y_out(stage_1_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({114906207, 95956458, 93815079, 119248786, 244981517, 25402945, 164849679, 253446904,
              182759226, 65939487, 218411001, 105651679, 13136617, 86425411, 248430418, 104273059,
              48258409, 32326785, 86611832, 248049881, 220409117, 60951044, 98839404, 128923754,
              50041017, 51590619, 71466452, 81879124, 6839312, 50250252, 70993112, 202017141,
              77785137, 166705511, 159555178, 176106545, 168682489, 99151986, 45900567, 135965343,
              95745785, 196552678, 266184237, 36678208, 124689641, 250979164, 196076822, 242448751,
              142932928, 232700332, 26885190, 157159811, 187973069, 49412866, 195777196, 24169593,
              242906033, 123556687, 258128862, 66398989, 60114085, 79759830, 203861878, 47380903}))
  stage_1_butterfly_19 (
    .x_in(stage_0_per_out[38]),
    .y_in(stage_0_per_out[39]),
    .x_out(stage_1_per_in[38]),
    .y_out(stage_1_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({236173805, 218922070, 59945410, 88068083, 184394225, 224193580, 73580010, 38581987,
              38792404, 22320040, 216197112, 213462715, 114462613, 232970901, 264463333, 143364478,
              127281316, 167753662, 212643172, 182920379, 48499686, 145595829, 67780496, 120068412,
              79121294, 122372515, 4519531, 126673466, 233112987, 267701123, 118263349, 83665434,
              12994463, 106279827, 221333762, 261080375, 252329804, 115935405, 205553550, 237391515,
              154194427, 153619107, 246502592, 248921617, 103784724, 96644160, 257122505, 54591848,
              117082039, 205764394, 85879269, 230500375, 91384253, 166918201, 253166836, 58002164,
              222792306, 174707320, 19111856, 120623833, 233855133, 215876710, 74620568, 117068649}))
  stage_1_butterfly_20 (
    .x_in(stage_0_per_out[40]),
    .y_in(stage_0_per_out[41]),
    .x_out(stage_1_per_in[40]),
    .y_out(stage_1_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({236173805, 218922070, 59945410, 88068083, 184394225, 224193580, 73580010, 38581987,
              38792404, 22320040, 216197112, 213462715, 114462613, 232970901, 264463333, 143364478,
              127281316, 167753662, 212643172, 182920379, 48499686, 145595829, 67780496, 120068412,
              79121294, 122372515, 4519531, 126673466, 233112987, 267701123, 118263349, 83665434,
              12994463, 106279827, 221333762, 261080375, 252329804, 115935405, 205553550, 237391515,
              154194427, 153619107, 246502592, 248921617, 103784724, 96644160, 257122505, 54591848,
              117082039, 205764394, 85879269, 230500375, 91384253, 166918201, 253166836, 58002164,
              222792306, 174707320, 19111856, 120623833, 233855133, 215876710, 74620568, 117068649}))
  stage_1_butterfly_21 (
    .x_in(stage_0_per_out[42]),
    .y_in(stage_0_per_out[43]),
    .x_out(stage_1_per_in[42]),
    .y_out(stage_1_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({154634100, 158913333, 195704814, 176734838, 100279875, 145325214, 265093046, 11727916,
              64402402, 60782408, 22419281, 20002868, 130965208, 104683412, 239219986, 123982174,
              185120175, 254862428, 258398710, 86422302, 127264350, 95857789, 205236983, 63759475,
              105759020, 61255010, 65162419, 220487343, 199811874, 253117467, 3615863, 114664154,
              126437335, 78726832, 67459976, 175735543, 178639438, 104494180, 43817935, 7525756,
              219155874, 238828812, 209365645, 21397846, 87333346, 59853183, 95592544, 80415871,
              240329350, 243959994, 83440545, 44095704, 109752985, 213675734, 91771920, 83594289,
              252048491, 215932651, 23196483, 209775390, 45533578, 129973973, 153870377, 177655074}))
  stage_1_butterfly_22 (
    .x_in(stage_0_per_out[44]),
    .y_in(stage_0_per_out[45]),
    .x_out(stage_1_per_in[44]),
    .y_out(stage_1_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({154634100, 158913333, 195704814, 176734838, 100279875, 145325214, 265093046, 11727916,
              64402402, 60782408, 22419281, 20002868, 130965208, 104683412, 239219986, 123982174,
              185120175, 254862428, 258398710, 86422302, 127264350, 95857789, 205236983, 63759475,
              105759020, 61255010, 65162419, 220487343, 199811874, 253117467, 3615863, 114664154,
              126437335, 78726832, 67459976, 175735543, 178639438, 104494180, 43817935, 7525756,
              219155874, 238828812, 209365645, 21397846, 87333346, 59853183, 95592544, 80415871,
              240329350, 243959994, 83440545, 44095704, 109752985, 213675734, 91771920, 83594289,
              252048491, 215932651, 23196483, 209775390, 45533578, 129973973, 153870377, 177655074}))
  stage_1_butterfly_23 (
    .x_in(stage_0_per_out[46]),
    .y_in(stage_0_per_out[47]),
    .x_out(stage_1_per_in[46]),
    .y_out(stage_1_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({82346526, 125480758, 58372872, 128081279, 226865216, 196727396, 5284602, 133543242,
              30998042, 53716996, 182147827, 26713518, 1381761, 171508784, 57884406, 5028136,
              126629575, 267892175, 14425613, 50106553, 61366355, 14195884, 234435452, 73917671,
              189834774, 195995970, 193726599, 181264550, 224367752, 79252444, 260962587, 125264465,
              110001979, 264722248, 230614882, 232215778, 90833651, 18807047, 41031357, 79343207,
              223156719, 205816155, 102404987, 192939426, 93188095, 262718787, 95943159, 15406607,
              216344829, 116341913, 77043356, 148816114, 76840577, 145444168, 126638229, 258312618,
              175434645, 175360485, 228233519, 85861280, 21699914, 158406994, 149817301, 146642358}))
  stage_1_butterfly_24 (
    .x_in(stage_0_per_out[48]),
    .y_in(stage_0_per_out[49]),
    .x_out(stage_1_per_in[48]),
    .y_out(stage_1_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({82346526, 125480758, 58372872, 128081279, 226865216, 196727396, 5284602, 133543242,
              30998042, 53716996, 182147827, 26713518, 1381761, 171508784, 57884406, 5028136,
              126629575, 267892175, 14425613, 50106553, 61366355, 14195884, 234435452, 73917671,
              189834774, 195995970, 193726599, 181264550, 224367752, 79252444, 260962587, 125264465,
              110001979, 264722248, 230614882, 232215778, 90833651, 18807047, 41031357, 79343207,
              223156719, 205816155, 102404987, 192939426, 93188095, 262718787, 95943159, 15406607,
              216344829, 116341913, 77043356, 148816114, 76840577, 145444168, 126638229, 258312618,
              175434645, 175360485, 228233519, 85861280, 21699914, 158406994, 149817301, 146642358}))
  stage_1_butterfly_25 (
    .x_in(stage_0_per_out[50]),
    .y_in(stage_0_per_out[51]),
    .x_out(stage_1_per_in[50]),
    .y_out(stage_1_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({124972666, 59278718, 35010964, 48487396, 144113751, 8772869, 146661492, 34093582,
              248813222, 140980229, 209335538, 264638858, 64059298, 187469377, 95362545, 70333973,
              12562435, 100306740, 121954140, 202839194, 133033169, 178750844, 176649880, 132216843,
              200991325, 203006324, 191064173, 226857524, 11713205, 6515518, 24417340, 214119665,
              50422568, 22483780, 152117270, 52952054, 209487240, 119598304, 140766862, 176646986,
              199654780, 27342032, 237702991, 80711179, 53666796, 114157546, 200880844, 184171973,
              54194127, 104225870, 53103748, 85943438, 85925921, 146917464, 39159482, 239243318,
              82994670, 24889364, 151554022, 165873702, 131606898, 71397785, 185196127, 159375180}))
  stage_1_butterfly_26 (
    .x_in(stage_0_per_out[52]),
    .y_in(stage_0_per_out[53]),
    .x_out(stage_1_per_in[52]),
    .y_out(stage_1_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({124972666, 59278718, 35010964, 48487396, 144113751, 8772869, 146661492, 34093582,
              248813222, 140980229, 209335538, 264638858, 64059298, 187469377, 95362545, 70333973,
              12562435, 100306740, 121954140, 202839194, 133033169, 178750844, 176649880, 132216843,
              200991325, 203006324, 191064173, 226857524, 11713205, 6515518, 24417340, 214119665,
              50422568, 22483780, 152117270, 52952054, 209487240, 119598304, 140766862, 176646986,
              199654780, 27342032, 237702991, 80711179, 53666796, 114157546, 200880844, 184171973,
              54194127, 104225870, 53103748, 85943438, 85925921, 146917464, 39159482, 239243318,
              82994670, 24889364, 151554022, 165873702, 131606898, 71397785, 185196127, 159375180}))
  stage_1_butterfly_27 (
    .x_in(stage_0_per_out[54]),
    .y_in(stage_0_per_out[55]),
    .x_out(stage_1_per_in[54]),
    .y_out(stage_1_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({259902883, 64064097, 32769539, 136417444, 253791818, 157208225, 90415400, 182812696,
              141049304, 144089543, 201671086, 81774581, 69255389, 256522921, 148688834, 212200386,
              5071752, 50115805, 18362334, 96014882, 134836604, 223616593, 239800333, 241368847,
              94872102, 38129962, 77506253, 221869909, 124878920, 119697484, 163120146, 217885801,
              96098889, 259065776, 70871651, 41460117, 242696977, 25013575, 95276657, 71010071,
              203277373, 62424622, 28990836, 18485653, 16822583, 255875272, 122635188, 155632772,
              185121114, 134337294, 225384963, 139206238, 148548934, 176530780, 41573703, 127930513,
              231508432, 73886338, 94729012, 52942312, 189935724, 75752194, 243900215, 4980542}))
  stage_1_butterfly_28 (
    .x_in(stage_0_per_out[56]),
    .y_in(stage_0_per_out[57]),
    .x_out(stage_1_per_in[56]),
    .y_out(stage_1_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({259902883, 64064097, 32769539, 136417444, 253791818, 157208225, 90415400, 182812696,
              141049304, 144089543, 201671086, 81774581, 69255389, 256522921, 148688834, 212200386,
              5071752, 50115805, 18362334, 96014882, 134836604, 223616593, 239800333, 241368847,
              94872102, 38129962, 77506253, 221869909, 124878920, 119697484, 163120146, 217885801,
              96098889, 259065776, 70871651, 41460117, 242696977, 25013575, 95276657, 71010071,
              203277373, 62424622, 28990836, 18485653, 16822583, 255875272, 122635188, 155632772,
              185121114, 134337294, 225384963, 139206238, 148548934, 176530780, 41573703, 127930513,
              231508432, 73886338, 94729012, 52942312, 189935724, 75752194, 243900215, 4980542}))
  stage_1_butterfly_29 (
    .x_in(stage_0_per_out[58]),
    .y_in(stage_0_per_out[59]),
    .x_out(stage_1_per_in[58]),
    .y_out(stage_1_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({127717239, 135644103, 6456449, 157158700, 172630653, 51299486, 217483488, 254780782,
              137520333, 50213981, 139730465, 108532653, 248206642, 34242638, 22116392, 134518349,
              259334239, 152505970, 13394971, 187892585, 112174110, 254241553, 179888950, 256890018,
              16703359, 35688570, 197641184, 153805373, 143389876, 258225039, 74661667, 50021352,
              75588758, 209423491, 4184358, 179675005, 33161823, 31515852, 107466416, 244217621,
              14369566, 27456585, 243789725, 94477870, 133797547, 207692352, 38723858, 12048336,
              227177249, 48893661, 215351473, 102888853, 55952036, 157311612, 192111834, 116226,
              186728485, 187345691, 153057061, 106441080, 170437415, 126420356, 6554463, 101380813}))
  stage_1_butterfly_30 (
    .x_in(stage_0_per_out[60]),
    .y_in(stage_0_per_out[61]),
    .x_out(stage_1_per_in[60]),
    .y_out(stage_1_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({127717239, 135644103, 6456449, 157158700, 172630653, 51299486, 217483488, 254780782,
              137520333, 50213981, 139730465, 108532653, 248206642, 34242638, 22116392, 134518349,
              259334239, 152505970, 13394971, 187892585, 112174110, 254241553, 179888950, 256890018,
              16703359, 35688570, 197641184, 153805373, 143389876, 258225039, 74661667, 50021352,
              75588758, 209423491, 4184358, 179675005, 33161823, 31515852, 107466416, 244217621,
              14369566, 27456585, 243789725, 94477870, 133797547, 207692352, 38723858, 12048336,
              227177249, 48893661, 215351473, 102888853, 55952036, 157311612, 192111834, 116226,
              186728485, 187345691, 153057061, 106441080, 170437415, 126420356, 6554463, 101380813}))
  stage_1_butterfly_31 (
    .x_in(stage_0_per_out[62]),
    .y_in(stage_0_per_out[63]),
    .x_out(stage_1_per_in[62]),
    .y_out(stage_1_per_in[63]),
    .clk(clk),
    .rst(rst)
  );




  
  // TODO(Yang): stage 1 -> stage 2 permutation
  // FIXME: ignore butterfly units for now.
  stage_1_permutation #(
    .DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    .INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_1_2_per (
    .inData_0(stage_1_per_in[0]),
    .inData_1(stage_1_per_in[1]),
    .inData_2(stage_1_per_in[2]),
    .inData_3(stage_1_per_in[3]),
    .inData_4(stage_1_per_in[4]),
    .inData_5(stage_1_per_in[5]),
    .inData_6(stage_1_per_in[6]),
    .inData_7(stage_1_per_in[7]),
    .inData_8(stage_1_per_in[8]),
    .inData_9(stage_1_per_in[9]),
    .inData_10(stage_1_per_in[10]),
    .inData_11(stage_1_per_in[11]),
    .inData_12(stage_1_per_in[12]),
    .inData_13(stage_1_per_in[13]),
    .inData_14(stage_1_per_in[14]),
    .inData_15(stage_1_per_in[15]),
    .inData_16(stage_1_per_in[16]),
    .inData_17(stage_1_per_in[17]),
    .inData_18(stage_1_per_in[18]),
    .inData_19(stage_1_per_in[19]),
    .inData_20(stage_1_per_in[20]),
    .inData_21(stage_1_per_in[21]),
    .inData_22(stage_1_per_in[22]),
    .inData_23(stage_1_per_in[23]),
    .inData_24(stage_1_per_in[24]),
    .inData_25(stage_1_per_in[25]),
    .inData_26(stage_1_per_in[26]),
    .inData_27(stage_1_per_in[27]),
    .inData_28(stage_1_per_in[28]),
    .inData_29(stage_1_per_in[29]),
    .inData_30(stage_1_per_in[30]),
    .inData_31(stage_1_per_in[31]),
    .inData_32(stage_1_per_in[32]),
    .inData_33(stage_1_per_in[33]),
    .inData_34(stage_1_per_in[34]),
    .inData_35(stage_1_per_in[35]),
    .inData_36(stage_1_per_in[36]),
    .inData_37(stage_1_per_in[37]),
    .inData_38(stage_1_per_in[38]),
    .inData_39(stage_1_per_in[39]),
    .inData_40(stage_1_per_in[40]),
    .inData_41(stage_1_per_in[41]),
    .inData_42(stage_1_per_in[42]),
    .inData_43(stage_1_per_in[43]),
    .inData_44(stage_1_per_in[44]),
    .inData_45(stage_1_per_in[45]),
    .inData_46(stage_1_per_in[46]),
    .inData_47(stage_1_per_in[47]),
    .inData_48(stage_1_per_in[48]),
    .inData_49(stage_1_per_in[49]),
    .inData_50(stage_1_per_in[50]),
    .inData_51(stage_1_per_in[51]),
    .inData_52(stage_1_per_in[52]),
    .inData_53(stage_1_per_in[53]),
    .inData_54(stage_1_per_in[54]),
    .inData_55(stage_1_per_in[55]),
    .inData_56(stage_1_per_in[56]),
    .inData_57(stage_1_per_in[57]),
    .inData_58(stage_1_per_in[58]),
    .inData_59(stage_1_per_in[59]),
    .inData_60(stage_1_per_in[60]),
    .inData_61(stage_1_per_in[61]),
    .inData_62(stage_1_per_in[62]),
    .inData_63(stage_1_per_in[63]),
    .outData_0(stage_1_per_out[0]),
    .outData_1(stage_1_per_out[1]),
    .outData_2(stage_1_per_out[2]),
    .outData_3(stage_1_per_out[3]),
    .outData_4(stage_1_per_out[4]),
    .outData_5(stage_1_per_out[5]),
    .outData_6(stage_1_per_out[6]),
    .outData_7(stage_1_per_out[7]),
    .outData_8(stage_1_per_out[8]),
    .outData_9(stage_1_per_out[9]),
    .outData_10(stage_1_per_out[10]),
    .outData_11(stage_1_per_out[11]),
    .outData_12(stage_1_per_out[12]),
    .outData_13(stage_1_per_out[13]),
    .outData_14(stage_1_per_out[14]),
    .outData_15(stage_1_per_out[15]),
    .outData_16(stage_1_per_out[16]),
    .outData_17(stage_1_per_out[17]),
    .outData_18(stage_1_per_out[18]),
    .outData_19(stage_1_per_out[19]),
    .outData_20(stage_1_per_out[20]),
    .outData_21(stage_1_per_out[21]),
    .outData_22(stage_1_per_out[22]),
    .outData_23(stage_1_per_out[23]),
    .outData_24(stage_1_per_out[24]),
    .outData_25(stage_1_per_out[25]),
    .outData_26(stage_1_per_out[26]),
    .outData_27(stage_1_per_out[27]),
    .outData_28(stage_1_per_out[28]),
    .outData_29(stage_1_per_out[29]),
    .outData_30(stage_1_per_out[30]),
    .outData_31(stage_1_per_out[31]),
    .outData_32(stage_1_per_out[32]),
    .outData_33(stage_1_per_out[33]),
    .outData_34(stage_1_per_out[34]),
    .outData_35(stage_1_per_out[35]),
    .outData_36(stage_1_per_out[36]),
    .outData_37(stage_1_per_out[37]),
    .outData_38(stage_1_per_out[38]),
    .outData_39(stage_1_per_out[39]),
    .outData_40(stage_1_per_out[40]),
    .outData_41(stage_1_per_out[41]),
    .outData_42(stage_1_per_out[42]),
    .outData_43(stage_1_per_out[43]),
    .outData_44(stage_1_per_out[44]),
    .outData_45(stage_1_per_out[45]),
    .outData_46(stage_1_per_out[46]),
    .outData_47(stage_1_per_out[47]),
    .outData_48(stage_1_per_out[48]),
    .outData_49(stage_1_per_out[49]),
    .outData_50(stage_1_per_out[50]),
    .outData_51(stage_1_per_out[51]),
    .outData_52(stage_1_per_out[52]),
    .outData_53(stage_1_per_out[53]),
    .outData_54(stage_1_per_out[54]),
    .outData_55(stage_1_per_out[55]),
    .outData_56(stage_1_per_out[56]),
    .outData_57(stage_1_per_out[57]),
    .outData_58(stage_1_per_out[58]),
    .outData_59(stage_1_per_out[59]),
    .outData_60(stage_1_per_out[60]),
    .outData_61(stage_1_per_out[61]),
    .outData_62(stage_1_per_out[62]),
    .outData_63(stage_1_per_out[63]),
    .in_start(in_start[1]),
    .out_start(out_start[1]),
    .clk(clk),
    .rst(rst)
  );


  // TODO(Tian): stage 2 32 butterfly units
  butterfly #(
    .start(START_CYCLE[2]),
    .factors({187381670, 235273242, 120217110, 135902522, 54714468, 249576229, 142656304, 122969043,
              196018390, 206341936, 212112171, 81414740, 26068775, 141956852, 174191574, 209112367,
              27439037, 72369588, 189139684, 265348407, 58661398, 1855205, 128297265, 171206517,
              174612628, 226834391, 23442787, 77127228, 35629855, 43000087, 50083600, 246787643,
              233083676, 237125965, 24365404, 244423105, 173628384, 85740049, 63661975, 90687088,
              142941966, 167645260, 252714435, 145831337, 10646661, 206116619, 156195364, 191744986,
              250031819, 121730405, 183613005, 205856513, 206844979, 174028560, 78273516, 175598948,
              121414397, 4721397, 72509307, 146344523, 255478273, 62435894, 255463943, 193174373}))
  stage_2_butterfly_0 (
    .x_in(stage_1_per_out[0]),
    .y_in(stage_1_per_out[1]),
    .x_out(stage_2_per_in[0]),
    .y_out(stage_2_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({187381670, 235273242, 120217110, 135902522, 54714468, 249576229, 142656304, 122969043,
              196018390, 206341936, 212112171, 81414740, 26068775, 141956852, 174191574, 209112367,
              27439037, 72369588, 189139684, 265348407, 58661398, 1855205, 128297265, 171206517,
              174612628, 226834391, 23442787, 77127228, 35629855, 43000087, 50083600, 246787643,
              233083676, 237125965, 24365404, 244423105, 173628384, 85740049, 63661975, 90687088,
              142941966, 167645260, 252714435, 145831337, 10646661, 206116619, 156195364, 191744986,
              250031819, 121730405, 183613005, 205856513, 206844979, 174028560, 78273516, 175598948,
              121414397, 4721397, 72509307, 146344523, 255478273, 62435894, 255463943, 193174373}))
  stage_2_butterfly_1 (
    .x_in(stage_1_per_out[2]),
    .y_in(stage_1_per_out[3]),
    .x_out(stage_2_per_in[2]),
    .y_out(stage_2_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({187381670, 235273242, 120217110, 135902522, 54714468, 249576229, 142656304, 122969043,
              196018390, 206341936, 212112171, 81414740, 26068775, 141956852, 174191574, 209112367,
              27439037, 72369588, 189139684, 265348407, 58661398, 1855205, 128297265, 171206517,
              174612628, 226834391, 23442787, 77127228, 35629855, 43000087, 50083600, 246787643,
              233083676, 237125965, 24365404, 244423105, 173628384, 85740049, 63661975, 90687088,
              142941966, 167645260, 252714435, 145831337, 10646661, 206116619, 156195364, 191744986,
              250031819, 121730405, 183613005, 205856513, 206844979, 174028560, 78273516, 175598948,
              121414397, 4721397, 72509307, 146344523, 255478273, 62435894, 255463943, 193174373}))
  stage_2_butterfly_2 (
    .x_in(stage_1_per_out[4]),
    .y_in(stage_1_per_out[5]),
    .x_out(stage_2_per_in[4]),
    .y_out(stage_2_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({187381670, 235273242, 120217110, 135902522, 54714468, 249576229, 142656304, 122969043,
              196018390, 206341936, 212112171, 81414740, 26068775, 141956852, 174191574, 209112367,
              27439037, 72369588, 189139684, 265348407, 58661398, 1855205, 128297265, 171206517,
              174612628, 226834391, 23442787, 77127228, 35629855, 43000087, 50083600, 246787643,
              233083676, 237125965, 24365404, 244423105, 173628384, 85740049, 63661975, 90687088,
              142941966, 167645260, 252714435, 145831337, 10646661, 206116619, 156195364, 191744986,
              250031819, 121730405, 183613005, 205856513, 206844979, 174028560, 78273516, 175598948,
              121414397, 4721397, 72509307, 146344523, 255478273, 62435894, 255463943, 193174373}))
  stage_2_butterfly_3 (
    .x_in(stage_1_per_out[6]),
    .y_in(stage_1_per_out[7]),
    .x_out(stage_2_per_in[6]),
    .y_out(stage_2_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({222912429, 77536776, 248922055, 189601976, 38252193, 155363318, 157839041, 94792077,
              243009216, 65889055, 21649526, 164248031, 187208958, 212237706, 116527240, 261541195,
              189909138, 205242220, 190586128, 34052825, 224322272, 86359417, 130154791, 254842567,
              75993973, 169792793, 259621463, 146205579, 509728, 256834872, 190565686, 159538295,
              82779345, 250727821, 211982342, 243339369, 58491201, 56723699, 147903734, 224922683,
              128589211, 191250025, 165001005, 136179523, 267008435, 61322741, 147014646, 57946842,
              54690936, 100611174, 174163034, 56545684, 53284215, 148479452, 226025718, 161217010,
              156298941, 141267184, 73072346, 5739737, 186048173, 223481427, 112360014, 103896237}))
  stage_2_butterfly_4 (
    .x_in(stage_1_per_out[8]),
    .y_in(stage_1_per_out[9]),
    .x_out(stage_2_per_in[8]),
    .y_out(stage_2_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({222912429, 77536776, 248922055, 189601976, 38252193, 155363318, 157839041, 94792077,
              243009216, 65889055, 21649526, 164248031, 187208958, 212237706, 116527240, 261541195,
              189909138, 205242220, 190586128, 34052825, 224322272, 86359417, 130154791, 254842567,
              75993973, 169792793, 259621463, 146205579, 509728, 256834872, 190565686, 159538295,
              82779345, 250727821, 211982342, 243339369, 58491201, 56723699, 147903734, 224922683,
              128589211, 191250025, 165001005, 136179523, 267008435, 61322741, 147014646, 57946842,
              54690936, 100611174, 174163034, 56545684, 53284215, 148479452, 226025718, 161217010,
              156298941, 141267184, 73072346, 5739737, 186048173, 223481427, 112360014, 103896237}))
  stage_2_butterfly_5 (
    .x_in(stage_1_per_out[10]),
    .y_in(stage_1_per_out[11]),
    .x_out(stage_2_per_in[10]),
    .y_out(stage_2_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({222912429, 77536776, 248922055, 189601976, 38252193, 155363318, 157839041, 94792077,
              243009216, 65889055, 21649526, 164248031, 187208958, 212237706, 116527240, 261541195,
              189909138, 205242220, 190586128, 34052825, 224322272, 86359417, 130154791, 254842567,
              75993973, 169792793, 259621463, 146205579, 509728, 256834872, 190565686, 159538295,
              82779345, 250727821, 211982342, 243339369, 58491201, 56723699, 147903734, 224922683,
              128589211, 191250025, 165001005, 136179523, 267008435, 61322741, 147014646, 57946842,
              54690936, 100611174, 174163034, 56545684, 53284215, 148479452, 226025718, 161217010,
              156298941, 141267184, 73072346, 5739737, 186048173, 223481427, 112360014, 103896237}))
  stage_2_butterfly_6 (
    .x_in(stage_1_per_out[12]),
    .y_in(stage_1_per_out[13]),
    .x_out(stage_2_per_in[12]),
    .y_out(stage_2_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({222912429, 77536776, 248922055, 189601976, 38252193, 155363318, 157839041, 94792077,
              243009216, 65889055, 21649526, 164248031, 187208958, 212237706, 116527240, 261541195,
              189909138, 205242220, 190586128, 34052825, 224322272, 86359417, 130154791, 254842567,
              75993973, 169792793, 259621463, 146205579, 509728, 256834872, 190565686, 159538295,
              82779345, 250727821, 211982342, 243339369, 58491201, 56723699, 147903734, 224922683,
              128589211, 191250025, 165001005, 136179523, 267008435, 61322741, 147014646, 57946842,
              54690936, 100611174, 174163034, 56545684, 53284215, 148479452, 226025718, 161217010,
              156298941, 141267184, 73072346, 5739737, 186048173, 223481427, 112360014, 103896237}))
  stage_2_butterfly_7 (
    .x_in(stage_1_per_out[14]),
    .y_in(stage_1_per_out[15]),
    .x_out(stage_2_per_in[14]),
    .y_out(stage_2_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({224391994, 73481957, 29779638, 116513948, 217763430, 89028484, 107830842, 187106042,
              193911793, 207877484, 168470500, 58903295, 267506256, 12286825, 82483914, 77916555,
              231354349, 181167176, 133273987, 145351880, 149788353, 160204962, 6760936, 45355620,
              54916848, 129325164, 207530748, 259302720, 36492987, 51550886, 91458750, 110378476,
              202032572, 218380292, 69017626, 140358303, 139374293, 3260661, 268043824, 19058782,
              158314046, 190540901, 121608761, 222527593, 153237233, 60600589, 159491687, 202565947,
              19700796, 50174239, 8474832, 226759664, 81838336, 46197346, 148491526, 92902456,
              13228372, 78552959, 255552842, 159148996, 8836114, 76313029, 256519333, 24036023}))
  stage_2_butterfly_8 (
    .x_in(stage_1_per_out[16]),
    .y_in(stage_1_per_out[17]),
    .x_out(stage_2_per_in[16]),
    .y_out(stage_2_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({224391994, 73481957, 29779638, 116513948, 217763430, 89028484, 107830842, 187106042,
              193911793, 207877484, 168470500, 58903295, 267506256, 12286825, 82483914, 77916555,
              231354349, 181167176, 133273987, 145351880, 149788353, 160204962, 6760936, 45355620,
              54916848, 129325164, 207530748, 259302720, 36492987, 51550886, 91458750, 110378476,
              202032572, 218380292, 69017626, 140358303, 139374293, 3260661, 268043824, 19058782,
              158314046, 190540901, 121608761, 222527593, 153237233, 60600589, 159491687, 202565947,
              19700796, 50174239, 8474832, 226759664, 81838336, 46197346, 148491526, 92902456,
              13228372, 78552959, 255552842, 159148996, 8836114, 76313029, 256519333, 24036023}))
  stage_2_butterfly_9 (
    .x_in(stage_1_per_out[18]),
    .y_in(stage_1_per_out[19]),
    .x_out(stage_2_per_in[18]),
    .y_out(stage_2_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({224391994, 73481957, 29779638, 116513948, 217763430, 89028484, 107830842, 187106042,
              193911793, 207877484, 168470500, 58903295, 267506256, 12286825, 82483914, 77916555,
              231354349, 181167176, 133273987, 145351880, 149788353, 160204962, 6760936, 45355620,
              54916848, 129325164, 207530748, 259302720, 36492987, 51550886, 91458750, 110378476,
              202032572, 218380292, 69017626, 140358303, 139374293, 3260661, 268043824, 19058782,
              158314046, 190540901, 121608761, 222527593, 153237233, 60600589, 159491687, 202565947,
              19700796, 50174239, 8474832, 226759664, 81838336, 46197346, 148491526, 92902456,
              13228372, 78552959, 255552842, 159148996, 8836114, 76313029, 256519333, 24036023}))
  stage_2_butterfly_10 (
    .x_in(stage_1_per_out[20]),
    .y_in(stage_1_per_out[21]),
    .x_out(stage_2_per_in[20]),
    .y_out(stage_2_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({224391994, 73481957, 29779638, 116513948, 217763430, 89028484, 107830842, 187106042,
              193911793, 207877484, 168470500, 58903295, 267506256, 12286825, 82483914, 77916555,
              231354349, 181167176, 133273987, 145351880, 149788353, 160204962, 6760936, 45355620,
              54916848, 129325164, 207530748, 259302720, 36492987, 51550886, 91458750, 110378476,
              202032572, 218380292, 69017626, 140358303, 139374293, 3260661, 268043824, 19058782,
              158314046, 190540901, 121608761, 222527593, 153237233, 60600589, 159491687, 202565947,
              19700796, 50174239, 8474832, 226759664, 81838336, 46197346, 148491526, 92902456,
              13228372, 78552959, 255552842, 159148996, 8836114, 76313029, 256519333, 24036023}))
  stage_2_butterfly_11 (
    .x_in(stage_1_per_out[22]),
    .y_in(stage_1_per_out[23]),
    .x_out(stage_2_per_in[22]),
    .y_out(stage_2_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({134161265, 183700349, 165671105, 188535281, 184464011, 174391063, 218207344, 266378632,
              236272786, 150049787, 33594840, 189044804, 197065781, 175710456, 14882191, 104215821,
              114052864, 159987098, 129677075, 140210175, 189757297, 72677507, 159978713, 197425604,
              171198428, 92441360, 195152646, 58726750, 99543252, 236050384, 94436408, 153319834,
              36196902, 135921552, 160050812, 161607031, 20655050, 9793208, 145034434, 52844710,
              233967292, 69205492, 134796549, 187867192, 184560259, 164728317, 99012968, 243091016,
              243047656, 8650362, 54393228, 8259535, 94686133, 79336225, 195270185, 234786570,
              249947221, 123052007, 132747224, 261458154, 237395333, 129740611, 227454343, 2204580}))
  stage_2_butterfly_12 (
    .x_in(stage_1_per_out[24]),
    .y_in(stage_1_per_out[25]),
    .x_out(stage_2_per_in[24]),
    .y_out(stage_2_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({134161265, 183700349, 165671105, 188535281, 184464011, 174391063, 218207344, 266378632,
              236272786, 150049787, 33594840, 189044804, 197065781, 175710456, 14882191, 104215821,
              114052864, 159987098, 129677075, 140210175, 189757297, 72677507, 159978713, 197425604,
              171198428, 92441360, 195152646, 58726750, 99543252, 236050384, 94436408, 153319834,
              36196902, 135921552, 160050812, 161607031, 20655050, 9793208, 145034434, 52844710,
              233967292, 69205492, 134796549, 187867192, 184560259, 164728317, 99012968, 243091016,
              243047656, 8650362, 54393228, 8259535, 94686133, 79336225, 195270185, 234786570,
              249947221, 123052007, 132747224, 261458154, 237395333, 129740611, 227454343, 2204580}))
  stage_2_butterfly_13 (
    .x_in(stage_1_per_out[26]),
    .y_in(stage_1_per_out[27]),
    .x_out(stage_2_per_in[26]),
    .y_out(stage_2_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({134161265, 183700349, 165671105, 188535281, 184464011, 174391063, 218207344, 266378632,
              236272786, 150049787, 33594840, 189044804, 197065781, 175710456, 14882191, 104215821,
              114052864, 159987098, 129677075, 140210175, 189757297, 72677507, 159978713, 197425604,
              171198428, 92441360, 195152646, 58726750, 99543252, 236050384, 94436408, 153319834,
              36196902, 135921552, 160050812, 161607031, 20655050, 9793208, 145034434, 52844710,
              233967292, 69205492, 134796549, 187867192, 184560259, 164728317, 99012968, 243091016,
              243047656, 8650362, 54393228, 8259535, 94686133, 79336225, 195270185, 234786570,
              249947221, 123052007, 132747224, 261458154, 237395333, 129740611, 227454343, 2204580}))
  stage_2_butterfly_14 (
    .x_in(stage_1_per_out[28]),
    .y_in(stage_1_per_out[29]),
    .x_out(stage_2_per_in[28]),
    .y_out(stage_2_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({134161265, 183700349, 165671105, 188535281, 184464011, 174391063, 218207344, 266378632,
              236272786, 150049787, 33594840, 189044804, 197065781, 175710456, 14882191, 104215821,
              114052864, 159987098, 129677075, 140210175, 189757297, 72677507, 159978713, 197425604,
              171198428, 92441360, 195152646, 58726750, 99543252, 236050384, 94436408, 153319834,
              36196902, 135921552, 160050812, 161607031, 20655050, 9793208, 145034434, 52844710,
              233967292, 69205492, 134796549, 187867192, 184560259, 164728317, 99012968, 243091016,
              243047656, 8650362, 54393228, 8259535, 94686133, 79336225, 195270185, 234786570,
              249947221, 123052007, 132747224, 261458154, 237395333, 129740611, 227454343, 2204580}))
  stage_2_butterfly_15 (
    .x_in(stage_1_per_out[30]),
    .y_in(stage_1_per_out[31]),
    .x_out(stage_2_per_in[30]),
    .y_out(stage_2_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({64830196, 266562472, 70325928, 232847226, 163197321, 83977288, 102034957, 144502563,
              31964447, 262112169, 251717800, 107503597, 9205704, 217359458, 85566308, 184177651,
              148108490, 172401093, 237616434, 5161923, 128052734, 22997488, 113049121, 252018541,
              261143222, 584543, 211201491, 183571221, 151857114, 198336839, 53025186, 66582189,
              74918627, 142807968, 83194655, 174290656, 31540722, 87492030, 167181901, 22383105,
              32160642, 46312994, 38415865, 238775640, 264974639, 248328138, 36213609, 250611881,
              156534179, 209698557, 148649408, 227453822, 42575603, 93513491, 263102666, 169092523,
              47531240, 258059551, 212425161, 139742686, 19817676, 131659168, 25652741, 113269084}))
  stage_2_butterfly_16 (
    .x_in(stage_1_per_out[32]),
    .y_in(stage_1_per_out[33]),
    .x_out(stage_2_per_in[32]),
    .y_out(stage_2_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({64830196, 266562472, 70325928, 232847226, 163197321, 83977288, 102034957, 144502563,
              31964447, 262112169, 251717800, 107503597, 9205704, 217359458, 85566308, 184177651,
              148108490, 172401093, 237616434, 5161923, 128052734, 22997488, 113049121, 252018541,
              261143222, 584543, 211201491, 183571221, 151857114, 198336839, 53025186, 66582189,
              74918627, 142807968, 83194655, 174290656, 31540722, 87492030, 167181901, 22383105,
              32160642, 46312994, 38415865, 238775640, 264974639, 248328138, 36213609, 250611881,
              156534179, 209698557, 148649408, 227453822, 42575603, 93513491, 263102666, 169092523,
              47531240, 258059551, 212425161, 139742686, 19817676, 131659168, 25652741, 113269084}))
  stage_2_butterfly_17 (
    .x_in(stage_1_per_out[34]),
    .y_in(stage_1_per_out[35]),
    .x_out(stage_2_per_in[34]),
    .y_out(stage_2_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({64830196, 266562472, 70325928, 232847226, 163197321, 83977288, 102034957, 144502563,
              31964447, 262112169, 251717800, 107503597, 9205704, 217359458, 85566308, 184177651,
              148108490, 172401093, 237616434, 5161923, 128052734, 22997488, 113049121, 252018541,
              261143222, 584543, 211201491, 183571221, 151857114, 198336839, 53025186, 66582189,
              74918627, 142807968, 83194655, 174290656, 31540722, 87492030, 167181901, 22383105,
              32160642, 46312994, 38415865, 238775640, 264974639, 248328138, 36213609, 250611881,
              156534179, 209698557, 148649408, 227453822, 42575603, 93513491, 263102666, 169092523,
              47531240, 258059551, 212425161, 139742686, 19817676, 131659168, 25652741, 113269084}))
  stage_2_butterfly_18 (
    .x_in(stage_1_per_out[36]),
    .y_in(stage_1_per_out[37]),
    .x_out(stage_2_per_in[36]),
    .y_out(stage_2_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({64830196, 266562472, 70325928, 232847226, 163197321, 83977288, 102034957, 144502563,
              31964447, 262112169, 251717800, 107503597, 9205704, 217359458, 85566308, 184177651,
              148108490, 172401093, 237616434, 5161923, 128052734, 22997488, 113049121, 252018541,
              261143222, 584543, 211201491, 183571221, 151857114, 198336839, 53025186, 66582189,
              74918627, 142807968, 83194655, 174290656, 31540722, 87492030, 167181901, 22383105,
              32160642, 46312994, 38415865, 238775640, 264974639, 248328138, 36213609, 250611881,
              156534179, 209698557, 148649408, 227453822, 42575603, 93513491, 263102666, 169092523,
              47531240, 258059551, 212425161, 139742686, 19817676, 131659168, 25652741, 113269084}))
  stage_2_butterfly_19 (
    .x_in(stage_1_per_out[38]),
    .y_in(stage_1_per_out[39]),
    .x_out(stage_2_per_in[38]),
    .y_out(stage_2_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({62456195, 65498827, 139101859, 181593250, 18205961, 73685379, 107513427, 133098101,
              90701762, 245041907, 228715598, 133952844, 122609533, 69412414, 37504237, 149904904,
              157649589, 265496406, 102785717, 55947412, 123720956, 134561032, 212728405, 131471427,
              163812077, 228572460, 257402730, 121970089, 29537138, 186476418, 248946430, 120318911,
              129694458, 149925004, 222087036, 236528116, 183590673, 210373784, 111532362, 53126225,
              12711531, 137060289, 162575967, 255737752, 86752434, 4457103, 153316076, 157386503,
              61348732, 23776027, 67784869, 212162524, 168674209, 203905228, 199055975, 50376784,
              5368199, 203598031, 37377133, 134804553, 127918992, 193897399, 143811089, 149423455}))
  stage_2_butterfly_20 (
    .x_in(stage_1_per_out[40]),
    .y_in(stage_1_per_out[41]),
    .x_out(stage_2_per_in[40]),
    .y_out(stage_2_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({62456195, 65498827, 139101859, 181593250, 18205961, 73685379, 107513427, 133098101,
              90701762, 245041907, 228715598, 133952844, 122609533, 69412414, 37504237, 149904904,
              157649589, 265496406, 102785717, 55947412, 123720956, 134561032, 212728405, 131471427,
              163812077, 228572460, 257402730, 121970089, 29537138, 186476418, 248946430, 120318911,
              129694458, 149925004, 222087036, 236528116, 183590673, 210373784, 111532362, 53126225,
              12711531, 137060289, 162575967, 255737752, 86752434, 4457103, 153316076, 157386503,
              61348732, 23776027, 67784869, 212162524, 168674209, 203905228, 199055975, 50376784,
              5368199, 203598031, 37377133, 134804553, 127918992, 193897399, 143811089, 149423455}))
  stage_2_butterfly_21 (
    .x_in(stage_1_per_out[42]),
    .y_in(stage_1_per_out[43]),
    .x_out(stage_2_per_in[42]),
    .y_out(stage_2_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({62456195, 65498827, 139101859, 181593250, 18205961, 73685379, 107513427, 133098101,
              90701762, 245041907, 228715598, 133952844, 122609533, 69412414, 37504237, 149904904,
              157649589, 265496406, 102785717, 55947412, 123720956, 134561032, 212728405, 131471427,
              163812077, 228572460, 257402730, 121970089, 29537138, 186476418, 248946430, 120318911,
              129694458, 149925004, 222087036, 236528116, 183590673, 210373784, 111532362, 53126225,
              12711531, 137060289, 162575967, 255737752, 86752434, 4457103, 153316076, 157386503,
              61348732, 23776027, 67784869, 212162524, 168674209, 203905228, 199055975, 50376784,
              5368199, 203598031, 37377133, 134804553, 127918992, 193897399, 143811089, 149423455}))
  stage_2_butterfly_22 (
    .x_in(stage_1_per_out[44]),
    .y_in(stage_1_per_out[45]),
    .x_out(stage_2_per_in[44]),
    .y_out(stage_2_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({62456195, 65498827, 139101859, 181593250, 18205961, 73685379, 107513427, 133098101,
              90701762, 245041907, 228715598, 133952844, 122609533, 69412414, 37504237, 149904904,
              157649589, 265496406, 102785717, 55947412, 123720956, 134561032, 212728405, 131471427,
              163812077, 228572460, 257402730, 121970089, 29537138, 186476418, 248946430, 120318911,
              129694458, 149925004, 222087036, 236528116, 183590673, 210373784, 111532362, 53126225,
              12711531, 137060289, 162575967, 255737752, 86752434, 4457103, 153316076, 157386503,
              61348732, 23776027, 67784869, 212162524, 168674209, 203905228, 199055975, 50376784,
              5368199, 203598031, 37377133, 134804553, 127918992, 193897399, 143811089, 149423455}))
  stage_2_butterfly_23 (
    .x_in(stage_1_per_out[46]),
    .y_in(stage_1_per_out[47]),
    .x_out(stage_2_per_in[46]),
    .y_out(stage_2_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({48885659, 98410858, 205681680, 16697663, 46120362, 163823140, 175949223, 56081948,
              233437339, 121712648, 127163336, 53432143, 79843127, 265883664, 90149574, 94856770,
              158914825, 126807666, 248133554, 23586243, 264322432, 123313741, 229032903, 232038388,
              7376627, 217846048, 4643973, 106743034, 120080647, 121145061, 98269185, 2487567,
              92379159, 6001670, 160048836, 55581691, 184522009, 170230234, 254234203, 180764097,
              100343421, 103503994, 195181845, 37498403, 66412546, 99996719, 126749676, 5445105,
              247452694, 62094530, 266777211, 219133933, 12551837, 55222727, 161345834, 183669067,
              255457916, 263649093, 59214954, 101579460, 110302060, 7301415, 135080569, 168342750}))
  stage_2_butterfly_24 (
    .x_in(stage_1_per_out[48]),
    .y_in(stage_1_per_out[49]),
    .x_out(stage_2_per_in[48]),
    .y_out(stage_2_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({48885659, 98410858, 205681680, 16697663, 46120362, 163823140, 175949223, 56081948,
              233437339, 121712648, 127163336, 53432143, 79843127, 265883664, 90149574, 94856770,
              158914825, 126807666, 248133554, 23586243, 264322432, 123313741, 229032903, 232038388,
              7376627, 217846048, 4643973, 106743034, 120080647, 121145061, 98269185, 2487567,
              92379159, 6001670, 160048836, 55581691, 184522009, 170230234, 254234203, 180764097,
              100343421, 103503994, 195181845, 37498403, 66412546, 99996719, 126749676, 5445105,
              247452694, 62094530, 266777211, 219133933, 12551837, 55222727, 161345834, 183669067,
              255457916, 263649093, 59214954, 101579460, 110302060, 7301415, 135080569, 168342750}))
  stage_2_butterfly_25 (
    .x_in(stage_1_per_out[50]),
    .y_in(stage_1_per_out[51]),
    .x_out(stage_2_per_in[50]),
    .y_out(stage_2_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({48885659, 98410858, 205681680, 16697663, 46120362, 163823140, 175949223, 56081948,
              233437339, 121712648, 127163336, 53432143, 79843127, 265883664, 90149574, 94856770,
              158914825, 126807666, 248133554, 23586243, 264322432, 123313741, 229032903, 232038388,
              7376627, 217846048, 4643973, 106743034, 120080647, 121145061, 98269185, 2487567,
              92379159, 6001670, 160048836, 55581691, 184522009, 170230234, 254234203, 180764097,
              100343421, 103503994, 195181845, 37498403, 66412546, 99996719, 126749676, 5445105,
              247452694, 62094530, 266777211, 219133933, 12551837, 55222727, 161345834, 183669067,
              255457916, 263649093, 59214954, 101579460, 110302060, 7301415, 135080569, 168342750}))
  stage_2_butterfly_26 (
    .x_in(stage_1_per_out[52]),
    .y_in(stage_1_per_out[53]),
    .x_out(stage_2_per_in[52]),
    .y_out(stage_2_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({48885659, 98410858, 205681680, 16697663, 46120362, 163823140, 175949223, 56081948,
              233437339, 121712648, 127163336, 53432143, 79843127, 265883664, 90149574, 94856770,
              158914825, 126807666, 248133554, 23586243, 264322432, 123313741, 229032903, 232038388,
              7376627, 217846048, 4643973, 106743034, 120080647, 121145061, 98269185, 2487567,
              92379159, 6001670, 160048836, 55581691, 184522009, 170230234, 254234203, 180764097,
              100343421, 103503994, 195181845, 37498403, 66412546, 99996719, 126749676, 5445105,
              247452694, 62094530, 266777211, 219133933, 12551837, 55222727, 161345834, 183669067,
              255457916, 263649093, 59214954, 101579460, 110302060, 7301415, 135080569, 168342750}))
  stage_2_butterfly_27 (
    .x_in(stage_1_per_out[54]),
    .y_in(stage_1_per_out[55]),
    .x_out(stage_2_per_in[54]),
    .y_out(stage_2_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({2017030, 217210388, 166139329, 17682401, 20118393, 60051251, 112756762, 107138937,
              95713937, 209744644, 224550271, 86350556, 67209795, 112825183, 248465751, 24347842,
              216531417, 62765404, 171841734, 19637177, 10943590, 81197166, 7280660, 244216061,
              267017218, 223473865, 105443909, 29901564, 154298223, 160429892, 247116469, 30998914,
              227628318, 102243739, 138513718, 21628090, 166586238, 226981541, 75689102, 95654178,
              195298807, 198352904, 266777383, 189248215, 265028258, 103189081, 151297332, 231749609,
              228243008, 58589536, 104290760, 74931497, 67241659, 255778637, 176972907, 178382895,
              116257755, 80381167, 27298769, 203850982, 122455193, 18433789, 208475153, 98445813}))
  stage_2_butterfly_28 (
    .x_in(stage_1_per_out[56]),
    .y_in(stage_1_per_out[57]),
    .x_out(stage_2_per_in[56]),
    .y_out(stage_2_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({2017030, 217210388, 166139329, 17682401, 20118393, 60051251, 112756762, 107138937,
              95713937, 209744644, 224550271, 86350556, 67209795, 112825183, 248465751, 24347842,
              216531417, 62765404, 171841734, 19637177, 10943590, 81197166, 7280660, 244216061,
              267017218, 223473865, 105443909, 29901564, 154298223, 160429892, 247116469, 30998914,
              227628318, 102243739, 138513718, 21628090, 166586238, 226981541, 75689102, 95654178,
              195298807, 198352904, 266777383, 189248215, 265028258, 103189081, 151297332, 231749609,
              228243008, 58589536, 104290760, 74931497, 67241659, 255778637, 176972907, 178382895,
              116257755, 80381167, 27298769, 203850982, 122455193, 18433789, 208475153, 98445813}))
  stage_2_butterfly_29 (
    .x_in(stage_1_per_out[58]),
    .y_in(stage_1_per_out[59]),
    .x_out(stage_2_per_in[58]),
    .y_out(stage_2_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({2017030, 217210388, 166139329, 17682401, 20118393, 60051251, 112756762, 107138937,
              95713937, 209744644, 224550271, 86350556, 67209795, 112825183, 248465751, 24347842,
              216531417, 62765404, 171841734, 19637177, 10943590, 81197166, 7280660, 244216061,
              267017218, 223473865, 105443909, 29901564, 154298223, 160429892, 247116469, 30998914,
              227628318, 102243739, 138513718, 21628090, 166586238, 226981541, 75689102, 95654178,
              195298807, 198352904, 266777383, 189248215, 265028258, 103189081, 151297332, 231749609,
              228243008, 58589536, 104290760, 74931497, 67241659, 255778637, 176972907, 178382895,
              116257755, 80381167, 27298769, 203850982, 122455193, 18433789, 208475153, 98445813}))
  stage_2_butterfly_30 (
    .x_in(stage_1_per_out[60]),
    .y_in(stage_1_per_out[61]),
    .x_out(stage_2_per_in[60]),
    .y_out(stage_2_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({2017030, 217210388, 166139329, 17682401, 20118393, 60051251, 112756762, 107138937,
              95713937, 209744644, 224550271, 86350556, 67209795, 112825183, 248465751, 24347842,
              216531417, 62765404, 171841734, 19637177, 10943590, 81197166, 7280660, 244216061,
              267017218, 223473865, 105443909, 29901564, 154298223, 160429892, 247116469, 30998914,
              227628318, 102243739, 138513718, 21628090, 166586238, 226981541, 75689102, 95654178,
              195298807, 198352904, 266777383, 189248215, 265028258, 103189081, 151297332, 231749609,
              228243008, 58589536, 104290760, 74931497, 67241659, 255778637, 176972907, 178382895,
              116257755, 80381167, 27298769, 203850982, 122455193, 18433789, 208475153, 98445813}))
  stage_2_butterfly_31 (
    .x_in(stage_1_per_out[62]),
    .y_in(stage_1_per_out[63]),
    .x_out(stage_2_per_in[62]),
    .y_out(stage_2_per_in[63]),
    .clk(clk),
    .rst(rst)
  );




  // TODO(Yang): stage 2 -> stage 3 permutation
  // FIXME: ignore butterfly units for now.
  stage_2_permutation #(
    .DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    .INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_2_3_per (
    .inData_0(stage_2_per_in[0]),
    .inData_1(stage_2_per_in[1]),
    .inData_2(stage_2_per_in[2]),
    .inData_3(stage_2_per_in[3]),
    .inData_4(stage_2_per_in[4]),
    .inData_5(stage_2_per_in[5]),
    .inData_6(stage_2_per_in[6]),
    .inData_7(stage_2_per_in[7]),
    .inData_8(stage_2_per_in[8]),
    .inData_9(stage_2_per_in[9]),
    .inData_10(stage_2_per_in[10]),
    .inData_11(stage_2_per_in[11]),
    .inData_12(stage_2_per_in[12]),
    .inData_13(stage_2_per_in[13]),
    .inData_14(stage_2_per_in[14]),
    .inData_15(stage_2_per_in[15]),
    .inData_16(stage_2_per_in[16]),
    .inData_17(stage_2_per_in[17]),
    .inData_18(stage_2_per_in[18]),
    .inData_19(stage_2_per_in[19]),
    .inData_20(stage_2_per_in[20]),
    .inData_21(stage_2_per_in[21]),
    .inData_22(stage_2_per_in[22]),
    .inData_23(stage_2_per_in[23]),
    .inData_24(stage_2_per_in[24]),
    .inData_25(stage_2_per_in[25]),
    .inData_26(stage_2_per_in[26]),
    .inData_27(stage_2_per_in[27]),
    .inData_28(stage_2_per_in[28]),
    .inData_29(stage_2_per_in[29]),
    .inData_30(stage_2_per_in[30]),
    .inData_31(stage_2_per_in[31]),
    .inData_32(stage_2_per_in[32]),
    .inData_33(stage_2_per_in[33]),
    .inData_34(stage_2_per_in[34]),
    .inData_35(stage_2_per_in[35]),
    .inData_36(stage_2_per_in[36]),
    .inData_37(stage_2_per_in[37]),
    .inData_38(stage_2_per_in[38]),
    .inData_39(stage_2_per_in[39]),
    .inData_40(stage_2_per_in[40]),
    .inData_41(stage_2_per_in[41]),
    .inData_42(stage_2_per_in[42]),
    .inData_43(stage_2_per_in[43]),
    .inData_44(stage_2_per_in[44]),
    .inData_45(stage_2_per_in[45]),
    .inData_46(stage_2_per_in[46]),
    .inData_47(stage_2_per_in[47]),
    .inData_48(stage_2_per_in[48]),
    .inData_49(stage_2_per_in[49]),
    .inData_50(stage_2_per_in[50]),
    .inData_51(stage_2_per_in[51]),
    .inData_52(stage_2_per_in[52]),
    .inData_53(stage_2_per_in[53]),
    .inData_54(stage_2_per_in[54]),
    .inData_55(stage_2_per_in[55]),
    .inData_56(stage_2_per_in[56]),
    .inData_57(stage_2_per_in[57]),
    .inData_58(stage_2_per_in[58]),
    .inData_59(stage_2_per_in[59]),
    .inData_60(stage_2_per_in[60]),
    .inData_61(stage_2_per_in[61]),
    .inData_62(stage_2_per_in[62]),
    .inData_63(stage_2_per_in[63]),
    .outData_0(stage_2_per_out[0]),
    .outData_1(stage_2_per_out[1]),
    .outData_2(stage_2_per_out[2]),
    .outData_3(stage_2_per_out[3]),
    .outData_4(stage_2_per_out[4]),
    .outData_5(stage_2_per_out[5]),
    .outData_6(stage_2_per_out[6]),
    .outData_7(stage_2_per_out[7]),
    .outData_8(stage_2_per_out[8]),
    .outData_9(stage_2_per_out[9]),
    .outData_10(stage_2_per_out[10]),
    .outData_11(stage_2_per_out[11]),
    .outData_12(stage_2_per_out[12]),
    .outData_13(stage_2_per_out[13]),
    .outData_14(stage_2_per_out[14]),
    .outData_15(stage_2_per_out[15]),
    .outData_16(stage_2_per_out[16]),
    .outData_17(stage_2_per_out[17]),
    .outData_18(stage_2_per_out[18]),
    .outData_19(stage_2_per_out[19]),
    .outData_20(stage_2_per_out[20]),
    .outData_21(stage_2_per_out[21]),
    .outData_22(stage_2_per_out[22]),
    .outData_23(stage_2_per_out[23]),
    .outData_24(stage_2_per_out[24]),
    .outData_25(stage_2_per_out[25]),
    .outData_26(stage_2_per_out[26]),
    .outData_27(stage_2_per_out[27]),
    .outData_28(stage_2_per_out[28]),
    .outData_29(stage_2_per_out[29]),
    .outData_30(stage_2_per_out[30]),
    .outData_31(stage_2_per_out[31]),
    .outData_32(stage_2_per_out[32]),
    .outData_33(stage_2_per_out[33]),
    .outData_34(stage_2_per_out[34]),
    .outData_35(stage_2_per_out[35]),
    .outData_36(stage_2_per_out[36]),
    .outData_37(stage_2_per_out[37]),
    .outData_38(stage_2_per_out[38]),
    .outData_39(stage_2_per_out[39]),
    .outData_40(stage_2_per_out[40]),
    .outData_41(stage_2_per_out[41]),
    .outData_42(stage_2_per_out[42]),
    .outData_43(stage_2_per_out[43]),
    .outData_44(stage_2_per_out[44]),
    .outData_45(stage_2_per_out[45]),
    .outData_46(stage_2_per_out[46]),
    .outData_47(stage_2_per_out[47]),
    .outData_48(stage_2_per_out[48]),
    .outData_49(stage_2_per_out[49]),
    .outData_50(stage_2_per_out[50]),
    .outData_51(stage_2_per_out[51]),
    .outData_52(stage_2_per_out[52]),
    .outData_53(stage_2_per_out[53]),
    .outData_54(stage_2_per_out[54]),
    .outData_55(stage_2_per_out[55]),
    .outData_56(stage_2_per_out[56]),
    .outData_57(stage_2_per_out[57]),
    .outData_58(stage_2_per_out[58]),
    .outData_59(stage_2_per_out[59]),
    .outData_60(stage_2_per_out[60]),
    .outData_61(stage_2_per_out[61]),
    .outData_62(stage_2_per_out[62]),
    .outData_63(stage_2_per_out[63]),
    .in_start(in_start[2]),
    .out_start(out_start[2]),
    .clk(clk),
    .rst(rst)
  );

  // TODO(Tian): stage 3 32 butterfly units
  butterfly #(
    .start(START_CYCLE[3]),
    .factors({135618975, 219738759, 141849606, 28242170, 98889920, 132483080, 134877507, 216395023,
              64884498, 42719459, 186863562, 168676526, 224068691, 212275822, 100123291, 190319963,
              209658551, 176209504, 99392088, 138879618, 258527796, 209725121, 85252512, 66242139,
              65324949, 49057739, 95282463, 262464837, 227819465, 183029478, 20857483, 80505160,
              198785423, 202059197, 1562592, 101414187, 219083512, 200399539, 194276347, 7460524,
              251898247, 34971158, 44144526, 103234978, 255286072, 206795535, 170930026, 171051327,
              224794776, 218231468, 176665584, 143969870, 202776751, 143779572, 246630386, 211426643,
              165872957, 247253507, 172508742, 242302870, 73698550, 25853611, 208297913, 36946189}))
  stage_3_butterfly_0 (
    .x_in(stage_2_per_out[0]),
    .y_in(stage_2_per_out[1]),
    .x_out(stage_3_per_in[0]),
    .y_out(stage_3_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({135618975, 219738759, 141849606, 28242170, 98889920, 132483080, 134877507, 216395023,
              64884498, 42719459, 186863562, 168676526, 224068691, 212275822, 100123291, 190319963,
              209658551, 176209504, 99392088, 138879618, 258527796, 209725121, 85252512, 66242139,
              65324949, 49057739, 95282463, 262464837, 227819465, 183029478, 20857483, 80505160,
              198785423, 202059197, 1562592, 101414187, 219083512, 200399539, 194276347, 7460524,
              251898247, 34971158, 44144526, 103234978, 255286072, 206795535, 170930026, 171051327,
              224794776, 218231468, 176665584, 143969870, 202776751, 143779572, 246630386, 211426643,
              165872957, 247253507, 172508742, 242302870, 73698550, 25853611, 208297913, 36946189}))
  stage_3_butterfly_1 (
    .x_in(stage_2_per_out[2]),
    .y_in(stage_2_per_out[3]),
    .x_out(stage_3_per_in[2]),
    .y_out(stage_3_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({135618975, 219738759, 141849606, 28242170, 98889920, 132483080, 134877507, 216395023,
              64884498, 42719459, 186863562, 168676526, 224068691, 212275822, 100123291, 190319963,
              209658551, 176209504, 99392088, 138879618, 258527796, 209725121, 85252512, 66242139,
              65324949, 49057739, 95282463, 262464837, 227819465, 183029478, 20857483, 80505160,
              198785423, 202059197, 1562592, 101414187, 219083512, 200399539, 194276347, 7460524,
              251898247, 34971158, 44144526, 103234978, 255286072, 206795535, 170930026, 171051327,
              224794776, 218231468, 176665584, 143969870, 202776751, 143779572, 246630386, 211426643,
              165872957, 247253507, 172508742, 242302870, 73698550, 25853611, 208297913, 36946189}))
  stage_3_butterfly_2 (
    .x_in(stage_2_per_out[4]),
    .y_in(stage_2_per_out[5]),
    .x_out(stage_3_per_in[4]),
    .y_out(stage_3_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({135618975, 219738759, 141849606, 28242170, 98889920, 132483080, 134877507, 216395023,
              64884498, 42719459, 186863562, 168676526, 224068691, 212275822, 100123291, 190319963,
              209658551, 176209504, 99392088, 138879618, 258527796, 209725121, 85252512, 66242139,
              65324949, 49057739, 95282463, 262464837, 227819465, 183029478, 20857483, 80505160,
              198785423, 202059197, 1562592, 101414187, 219083512, 200399539, 194276347, 7460524,
              251898247, 34971158, 44144526, 103234978, 255286072, 206795535, 170930026, 171051327,
              224794776, 218231468, 176665584, 143969870, 202776751, 143779572, 246630386, 211426643,
              165872957, 247253507, 172508742, 242302870, 73698550, 25853611, 208297913, 36946189}))
  stage_3_butterfly_3 (
    .x_in(stage_2_per_out[6]),
    .y_in(stage_2_per_out[7]),
    .x_out(stage_3_per_in[6]),
    .y_out(stage_3_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({135618975, 219738759, 141849606, 28242170, 98889920, 132483080, 134877507, 216395023,
              64884498, 42719459, 186863562, 168676526, 224068691, 212275822, 100123291, 190319963,
              209658551, 176209504, 99392088, 138879618, 258527796, 209725121, 85252512, 66242139,
              65324949, 49057739, 95282463, 262464837, 227819465, 183029478, 20857483, 80505160,
              198785423, 202059197, 1562592, 101414187, 219083512, 200399539, 194276347, 7460524,
              251898247, 34971158, 44144526, 103234978, 255286072, 206795535, 170930026, 171051327,
              224794776, 218231468, 176665584, 143969870, 202776751, 143779572, 246630386, 211426643,
              165872957, 247253507, 172508742, 242302870, 73698550, 25853611, 208297913, 36946189}))
  stage_3_butterfly_4 (
    .x_in(stage_2_per_out[8]),
    .y_in(stage_2_per_out[9]),
    .x_out(stage_3_per_in[8]),
    .y_out(stage_3_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({135618975, 219738759, 141849606, 28242170, 98889920, 132483080, 134877507, 216395023,
              64884498, 42719459, 186863562, 168676526, 224068691, 212275822, 100123291, 190319963,
              209658551, 176209504, 99392088, 138879618, 258527796, 209725121, 85252512, 66242139,
              65324949, 49057739, 95282463, 262464837, 227819465, 183029478, 20857483, 80505160,
              198785423, 202059197, 1562592, 101414187, 219083512, 200399539, 194276347, 7460524,
              251898247, 34971158, 44144526, 103234978, 255286072, 206795535, 170930026, 171051327,
              224794776, 218231468, 176665584, 143969870, 202776751, 143779572, 246630386, 211426643,
              165872957, 247253507, 172508742, 242302870, 73698550, 25853611, 208297913, 36946189}))
  stage_3_butterfly_5 (
    .x_in(stage_2_per_out[10]),
    .y_in(stage_2_per_out[11]),
    .x_out(stage_3_per_in[10]),
    .y_out(stage_3_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({135618975, 219738759, 141849606, 28242170, 98889920, 132483080, 134877507, 216395023,
              64884498, 42719459, 186863562, 168676526, 224068691, 212275822, 100123291, 190319963,
              209658551, 176209504, 99392088, 138879618, 258527796, 209725121, 85252512, 66242139,
              65324949, 49057739, 95282463, 262464837, 227819465, 183029478, 20857483, 80505160,
              198785423, 202059197, 1562592, 101414187, 219083512, 200399539, 194276347, 7460524,
              251898247, 34971158, 44144526, 103234978, 255286072, 206795535, 170930026, 171051327,
              224794776, 218231468, 176665584, 143969870, 202776751, 143779572, 246630386, 211426643,
              165872957, 247253507, 172508742, 242302870, 73698550, 25853611, 208297913, 36946189}))
  stage_3_butterfly_6 (
    .x_in(stage_2_per_out[12]),
    .y_in(stage_2_per_out[13]),
    .x_out(stage_3_per_in[12]),
    .y_out(stage_3_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({135618975, 219738759, 141849606, 28242170, 98889920, 132483080, 134877507, 216395023,
              64884498, 42719459, 186863562, 168676526, 224068691, 212275822, 100123291, 190319963,
              209658551, 176209504, 99392088, 138879618, 258527796, 209725121, 85252512, 66242139,
              65324949, 49057739, 95282463, 262464837, 227819465, 183029478, 20857483, 80505160,
              198785423, 202059197, 1562592, 101414187, 219083512, 200399539, 194276347, 7460524,
              251898247, 34971158, 44144526, 103234978, 255286072, 206795535, 170930026, 171051327,
              224794776, 218231468, 176665584, 143969870, 202776751, 143779572, 246630386, 211426643,
              165872957, 247253507, 172508742, 242302870, 73698550, 25853611, 208297913, 36946189}))
  stage_3_butterfly_7 (
    .x_in(stage_2_per_out[14]),
    .y_in(stage_2_per_out[15]),
    .x_out(stage_3_per_in[14]),
    .y_out(stage_3_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({42355602, 24688427, 45686070, 110403916, 78649100, 170284131, 17861009, 202071175,
              160254284, 224586596, 57574719, 181281889, 117221766, 205290416, 182702557, 65413984,
              136878682, 129576773, 5829490, 61644903, 61345534, 263077695, 148801771, 67321994,
              69773246, 196771169, 56155754, 82155735, 137065607, 155060883, 40158424, 207329882,
              54534442, 258226806, 249146534, 219898221, 61720173, 167366585, 64764693, 93469550,
              258559590, 68493159, 134269022, 63483304, 184644727, 225389748, 142306631, 95251863,
              220994759, 17231623, 8950678, 252241817, 225784463, 156366160, 61664240, 35918322,
              23892097, 35924353, 234350511, 6574921, 49504466, 119169851, 66505970, 6292910}))
  stage_3_butterfly_8 (
    .x_in(stage_2_per_out[16]),
    .y_in(stage_2_per_out[17]),
    .x_out(stage_3_per_in[16]),
    .y_out(stage_3_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({42355602, 24688427, 45686070, 110403916, 78649100, 170284131, 17861009, 202071175,
              160254284, 224586596, 57574719, 181281889, 117221766, 205290416, 182702557, 65413984,
              136878682, 129576773, 5829490, 61644903, 61345534, 263077695, 148801771, 67321994,
              69773246, 196771169, 56155754, 82155735, 137065607, 155060883, 40158424, 207329882,
              54534442, 258226806, 249146534, 219898221, 61720173, 167366585, 64764693, 93469550,
              258559590, 68493159, 134269022, 63483304, 184644727, 225389748, 142306631, 95251863,
              220994759, 17231623, 8950678, 252241817, 225784463, 156366160, 61664240, 35918322,
              23892097, 35924353, 234350511, 6574921, 49504466, 119169851, 66505970, 6292910}))
  stage_3_butterfly_9 (
    .x_in(stage_2_per_out[18]),
    .y_in(stage_2_per_out[19]),
    .x_out(stage_3_per_in[18]),
    .y_out(stage_3_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({42355602, 24688427, 45686070, 110403916, 78649100, 170284131, 17861009, 202071175,
              160254284, 224586596, 57574719, 181281889, 117221766, 205290416, 182702557, 65413984,
              136878682, 129576773, 5829490, 61644903, 61345534, 263077695, 148801771, 67321994,
              69773246, 196771169, 56155754, 82155735, 137065607, 155060883, 40158424, 207329882,
              54534442, 258226806, 249146534, 219898221, 61720173, 167366585, 64764693, 93469550,
              258559590, 68493159, 134269022, 63483304, 184644727, 225389748, 142306631, 95251863,
              220994759, 17231623, 8950678, 252241817, 225784463, 156366160, 61664240, 35918322,
              23892097, 35924353, 234350511, 6574921, 49504466, 119169851, 66505970, 6292910}))
  stage_3_butterfly_10 (
    .x_in(stage_2_per_out[20]),
    .y_in(stage_2_per_out[21]),
    .x_out(stage_3_per_in[20]),
    .y_out(stage_3_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({42355602, 24688427, 45686070, 110403916, 78649100, 170284131, 17861009, 202071175,
              160254284, 224586596, 57574719, 181281889, 117221766, 205290416, 182702557, 65413984,
              136878682, 129576773, 5829490, 61644903, 61345534, 263077695, 148801771, 67321994,
              69773246, 196771169, 56155754, 82155735, 137065607, 155060883, 40158424, 207329882,
              54534442, 258226806, 249146534, 219898221, 61720173, 167366585, 64764693, 93469550,
              258559590, 68493159, 134269022, 63483304, 184644727, 225389748, 142306631, 95251863,
              220994759, 17231623, 8950678, 252241817, 225784463, 156366160, 61664240, 35918322,
              23892097, 35924353, 234350511, 6574921, 49504466, 119169851, 66505970, 6292910}))
  stage_3_butterfly_11 (
    .x_in(stage_2_per_out[22]),
    .y_in(stage_2_per_out[23]),
    .x_out(stage_3_per_in[22]),
    .y_out(stage_3_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({42355602, 24688427, 45686070, 110403916, 78649100, 170284131, 17861009, 202071175,
              160254284, 224586596, 57574719, 181281889, 117221766, 205290416, 182702557, 65413984,
              136878682, 129576773, 5829490, 61644903, 61345534, 263077695, 148801771, 67321994,
              69773246, 196771169, 56155754, 82155735, 137065607, 155060883, 40158424, 207329882,
              54534442, 258226806, 249146534, 219898221, 61720173, 167366585, 64764693, 93469550,
              258559590, 68493159, 134269022, 63483304, 184644727, 225389748, 142306631, 95251863,
              220994759, 17231623, 8950678, 252241817, 225784463, 156366160, 61664240, 35918322,
              23892097, 35924353, 234350511, 6574921, 49504466, 119169851, 66505970, 6292910}))
  stage_3_butterfly_12 (
    .x_in(stage_2_per_out[24]),
    .y_in(stage_2_per_out[25]),
    .x_out(stage_3_per_in[24]),
    .y_out(stage_3_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({42355602, 24688427, 45686070, 110403916, 78649100, 170284131, 17861009, 202071175,
              160254284, 224586596, 57574719, 181281889, 117221766, 205290416, 182702557, 65413984,
              136878682, 129576773, 5829490, 61644903, 61345534, 263077695, 148801771, 67321994,
              69773246, 196771169, 56155754, 82155735, 137065607, 155060883, 40158424, 207329882,
              54534442, 258226806, 249146534, 219898221, 61720173, 167366585, 64764693, 93469550,
              258559590, 68493159, 134269022, 63483304, 184644727, 225389748, 142306631, 95251863,
              220994759, 17231623, 8950678, 252241817, 225784463, 156366160, 61664240, 35918322,
              23892097, 35924353, 234350511, 6574921, 49504466, 119169851, 66505970, 6292910}))
  stage_3_butterfly_13 (
    .x_in(stage_2_per_out[26]),
    .y_in(stage_2_per_out[27]),
    .x_out(stage_3_per_in[26]),
    .y_out(stage_3_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({42355602, 24688427, 45686070, 110403916, 78649100, 170284131, 17861009, 202071175,
              160254284, 224586596, 57574719, 181281889, 117221766, 205290416, 182702557, 65413984,
              136878682, 129576773, 5829490, 61644903, 61345534, 263077695, 148801771, 67321994,
              69773246, 196771169, 56155754, 82155735, 137065607, 155060883, 40158424, 207329882,
              54534442, 258226806, 249146534, 219898221, 61720173, 167366585, 64764693, 93469550,
              258559590, 68493159, 134269022, 63483304, 184644727, 225389748, 142306631, 95251863,
              220994759, 17231623, 8950678, 252241817, 225784463, 156366160, 61664240, 35918322,
              23892097, 35924353, 234350511, 6574921, 49504466, 119169851, 66505970, 6292910}))
  stage_3_butterfly_14 (
    .x_in(stage_2_per_out[28]),
    .y_in(stage_2_per_out[29]),
    .x_out(stage_3_per_in[28]),
    .y_out(stage_3_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({42355602, 24688427, 45686070, 110403916, 78649100, 170284131, 17861009, 202071175,
              160254284, 224586596, 57574719, 181281889, 117221766, 205290416, 182702557, 65413984,
              136878682, 129576773, 5829490, 61644903, 61345534, 263077695, 148801771, 67321994,
              69773246, 196771169, 56155754, 82155735, 137065607, 155060883, 40158424, 207329882,
              54534442, 258226806, 249146534, 219898221, 61720173, 167366585, 64764693, 93469550,
              258559590, 68493159, 134269022, 63483304, 184644727, 225389748, 142306631, 95251863,
              220994759, 17231623, 8950678, 252241817, 225784463, 156366160, 61664240, 35918322,
              23892097, 35924353, 234350511, 6574921, 49504466, 119169851, 66505970, 6292910}))
  stage_3_butterfly_15 (
    .x_in(stage_2_per_out[30]),
    .y_in(stage_2_per_out[31]),
    .x_out(stage_3_per_in[30]),
    .y_out(stage_3_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({98861208, 4839268, 12196542, 178386996, 232615475, 102915173, 201144768, 167911982,
              253800975, 263070789, 181295312, 131377029, 205961920, 82934386, 23606744, 76925614,
              79852752, 117274103, 32087335, 73081523, 141424302, 68267735, 172809179, 68559335,
              123440080, 55609416, 94612904, 190980049, 181468172, 243024363, 16985430, 195748297,
              233514072, 10720790, 185685569, 210770212, 172935357, 236109059, 44547301, 222861227,
              93740850, 225265815, 143102859, 256272276, 109902969, 47879495, 164638888, 177340471,
              87202272, 40718170, 57455860, 165350229, 150862394, 43194148, 161171966, 200749611,
              1613379, 256869432, 6010959, 209583375, 225291788, 139268485, 215146927, 257269778}))
  stage_3_butterfly_16 (
    .x_in(stage_2_per_out[32]),
    .y_in(stage_2_per_out[33]),
    .x_out(stage_3_per_in[32]),
    .y_out(stage_3_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({98861208, 4839268, 12196542, 178386996, 232615475, 102915173, 201144768, 167911982,
              253800975, 263070789, 181295312, 131377029, 205961920, 82934386, 23606744, 76925614,
              79852752, 117274103, 32087335, 73081523, 141424302, 68267735, 172809179, 68559335,
              123440080, 55609416, 94612904, 190980049, 181468172, 243024363, 16985430, 195748297,
              233514072, 10720790, 185685569, 210770212, 172935357, 236109059, 44547301, 222861227,
              93740850, 225265815, 143102859, 256272276, 109902969, 47879495, 164638888, 177340471,
              87202272, 40718170, 57455860, 165350229, 150862394, 43194148, 161171966, 200749611,
              1613379, 256869432, 6010959, 209583375, 225291788, 139268485, 215146927, 257269778}))
  stage_3_butterfly_17 (
    .x_in(stage_2_per_out[34]),
    .y_in(stage_2_per_out[35]),
    .x_out(stage_3_per_in[34]),
    .y_out(stage_3_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({98861208, 4839268, 12196542, 178386996, 232615475, 102915173, 201144768, 167911982,
              253800975, 263070789, 181295312, 131377029, 205961920, 82934386, 23606744, 76925614,
              79852752, 117274103, 32087335, 73081523, 141424302, 68267735, 172809179, 68559335,
              123440080, 55609416, 94612904, 190980049, 181468172, 243024363, 16985430, 195748297,
              233514072, 10720790, 185685569, 210770212, 172935357, 236109059, 44547301, 222861227,
              93740850, 225265815, 143102859, 256272276, 109902969, 47879495, 164638888, 177340471,
              87202272, 40718170, 57455860, 165350229, 150862394, 43194148, 161171966, 200749611,
              1613379, 256869432, 6010959, 209583375, 225291788, 139268485, 215146927, 257269778}))
  stage_3_butterfly_18 (
    .x_in(stage_2_per_out[36]),
    .y_in(stage_2_per_out[37]),
    .x_out(stage_3_per_in[36]),
    .y_out(stage_3_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({98861208, 4839268, 12196542, 178386996, 232615475, 102915173, 201144768, 167911982,
              253800975, 263070789, 181295312, 131377029, 205961920, 82934386, 23606744, 76925614,
              79852752, 117274103, 32087335, 73081523, 141424302, 68267735, 172809179, 68559335,
              123440080, 55609416, 94612904, 190980049, 181468172, 243024363, 16985430, 195748297,
              233514072, 10720790, 185685569, 210770212, 172935357, 236109059, 44547301, 222861227,
              93740850, 225265815, 143102859, 256272276, 109902969, 47879495, 164638888, 177340471,
              87202272, 40718170, 57455860, 165350229, 150862394, 43194148, 161171966, 200749611,
              1613379, 256869432, 6010959, 209583375, 225291788, 139268485, 215146927, 257269778}))
  stage_3_butterfly_19 (
    .x_in(stage_2_per_out[38]),
    .y_in(stage_2_per_out[39]),
    .x_out(stage_3_per_in[38]),
    .y_out(stage_3_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({98861208, 4839268, 12196542, 178386996, 232615475, 102915173, 201144768, 167911982,
              253800975, 263070789, 181295312, 131377029, 205961920, 82934386, 23606744, 76925614,
              79852752, 117274103, 32087335, 73081523, 141424302, 68267735, 172809179, 68559335,
              123440080, 55609416, 94612904, 190980049, 181468172, 243024363, 16985430, 195748297,
              233514072, 10720790, 185685569, 210770212, 172935357, 236109059, 44547301, 222861227,
              93740850, 225265815, 143102859, 256272276, 109902969, 47879495, 164638888, 177340471,
              87202272, 40718170, 57455860, 165350229, 150862394, 43194148, 161171966, 200749611,
              1613379, 256869432, 6010959, 209583375, 225291788, 139268485, 215146927, 257269778}))
  stage_3_butterfly_20 (
    .x_in(stage_2_per_out[40]),
    .y_in(stage_2_per_out[41]),
    .x_out(stage_3_per_in[40]),
    .y_out(stage_3_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({98861208, 4839268, 12196542, 178386996, 232615475, 102915173, 201144768, 167911982,
              253800975, 263070789, 181295312, 131377029, 205961920, 82934386, 23606744, 76925614,
              79852752, 117274103, 32087335, 73081523, 141424302, 68267735, 172809179, 68559335,
              123440080, 55609416, 94612904, 190980049, 181468172, 243024363, 16985430, 195748297,
              233514072, 10720790, 185685569, 210770212, 172935357, 236109059, 44547301, 222861227,
              93740850, 225265815, 143102859, 256272276, 109902969, 47879495, 164638888, 177340471,
              87202272, 40718170, 57455860, 165350229, 150862394, 43194148, 161171966, 200749611,
              1613379, 256869432, 6010959, 209583375, 225291788, 139268485, 215146927, 257269778}))
  stage_3_butterfly_21 (
    .x_in(stage_2_per_out[42]),
    .y_in(stage_2_per_out[43]),
    .x_out(stage_3_per_in[42]),
    .y_out(stage_3_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({98861208, 4839268, 12196542, 178386996, 232615475, 102915173, 201144768, 167911982,
              253800975, 263070789, 181295312, 131377029, 205961920, 82934386, 23606744, 76925614,
              79852752, 117274103, 32087335, 73081523, 141424302, 68267735, 172809179, 68559335,
              123440080, 55609416, 94612904, 190980049, 181468172, 243024363, 16985430, 195748297,
              233514072, 10720790, 185685569, 210770212, 172935357, 236109059, 44547301, 222861227,
              93740850, 225265815, 143102859, 256272276, 109902969, 47879495, 164638888, 177340471,
              87202272, 40718170, 57455860, 165350229, 150862394, 43194148, 161171966, 200749611,
              1613379, 256869432, 6010959, 209583375, 225291788, 139268485, 215146927, 257269778}))
  stage_3_butterfly_22 (
    .x_in(stage_2_per_out[44]),
    .y_in(stage_2_per_out[45]),
    .x_out(stage_3_per_in[44]),
    .y_out(stage_3_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({98861208, 4839268, 12196542, 178386996, 232615475, 102915173, 201144768, 167911982,
              253800975, 263070789, 181295312, 131377029, 205961920, 82934386, 23606744, 76925614,
              79852752, 117274103, 32087335, 73081523, 141424302, 68267735, 172809179, 68559335,
              123440080, 55609416, 94612904, 190980049, 181468172, 243024363, 16985430, 195748297,
              233514072, 10720790, 185685569, 210770212, 172935357, 236109059, 44547301, 222861227,
              93740850, 225265815, 143102859, 256272276, 109902969, 47879495, 164638888, 177340471,
              87202272, 40718170, 57455860, 165350229, 150862394, 43194148, 161171966, 200749611,
              1613379, 256869432, 6010959, 209583375, 225291788, 139268485, 215146927, 257269778}))
  stage_3_butterfly_23 (
    .x_in(stage_2_per_out[46]),
    .y_in(stage_2_per_out[47]),
    .x_out(stage_3_per_in[46]),
    .y_out(stage_3_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({77981460, 233888407, 199633043, 23405380, 142181410, 169182486, 160841949, 254132077,
              8411857, 34256894, 100229847, 79136411, 75073484, 109479656, 13458851, 205525433,
              192832423, 60548134, 56246211, 140366124, 62117518, 210734246, 148390399, 149992379,
              209085090, 50986641, 10003248, 114486793, 241313184, 266671862, 25944135, 184310992,
              212802310, 237102043, 50222736, 131023241, 18298478, 229100654, 209886001, 196522490,
              145034471, 185138250, 186841927, 122332647, 160807241, 247289727, 258257144, 196328787,
              193915204, 154421517, 92650808, 238382196, 171362072, 171541778, 30930936, 61997323,
              158727274, 242025902, 226213489, 137672988, 244216783, 49675259, 158168844, 182691070}))
  stage_3_butterfly_24 (
    .x_in(stage_2_per_out[48]),
    .y_in(stage_2_per_out[49]),
    .x_out(stage_3_per_in[48]),
    .y_out(stage_3_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({77981460, 233888407, 199633043, 23405380, 142181410, 169182486, 160841949, 254132077,
              8411857, 34256894, 100229847, 79136411, 75073484, 109479656, 13458851, 205525433,
              192832423, 60548134, 56246211, 140366124, 62117518, 210734246, 148390399, 149992379,
              209085090, 50986641, 10003248, 114486793, 241313184, 266671862, 25944135, 184310992,
              212802310, 237102043, 50222736, 131023241, 18298478, 229100654, 209886001, 196522490,
              145034471, 185138250, 186841927, 122332647, 160807241, 247289727, 258257144, 196328787,
              193915204, 154421517, 92650808, 238382196, 171362072, 171541778, 30930936, 61997323,
              158727274, 242025902, 226213489, 137672988, 244216783, 49675259, 158168844, 182691070}))
  stage_3_butterfly_25 (
    .x_in(stage_2_per_out[50]),
    .y_in(stage_2_per_out[51]),
    .x_out(stage_3_per_in[50]),
    .y_out(stage_3_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({77981460, 233888407, 199633043, 23405380, 142181410, 169182486, 160841949, 254132077,
              8411857, 34256894, 100229847, 79136411, 75073484, 109479656, 13458851, 205525433,
              192832423, 60548134, 56246211, 140366124, 62117518, 210734246, 148390399, 149992379,
              209085090, 50986641, 10003248, 114486793, 241313184, 266671862, 25944135, 184310992,
              212802310, 237102043, 50222736, 131023241, 18298478, 229100654, 209886001, 196522490,
              145034471, 185138250, 186841927, 122332647, 160807241, 247289727, 258257144, 196328787,
              193915204, 154421517, 92650808, 238382196, 171362072, 171541778, 30930936, 61997323,
              158727274, 242025902, 226213489, 137672988, 244216783, 49675259, 158168844, 182691070}))
  stage_3_butterfly_26 (
    .x_in(stage_2_per_out[52]),
    .y_in(stage_2_per_out[53]),
    .x_out(stage_3_per_in[52]),
    .y_out(stage_3_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({77981460, 233888407, 199633043, 23405380, 142181410, 169182486, 160841949, 254132077,
              8411857, 34256894, 100229847, 79136411, 75073484, 109479656, 13458851, 205525433,
              192832423, 60548134, 56246211, 140366124, 62117518, 210734246, 148390399, 149992379,
              209085090, 50986641, 10003248, 114486793, 241313184, 266671862, 25944135, 184310992,
              212802310, 237102043, 50222736, 131023241, 18298478, 229100654, 209886001, 196522490,
              145034471, 185138250, 186841927, 122332647, 160807241, 247289727, 258257144, 196328787,
              193915204, 154421517, 92650808, 238382196, 171362072, 171541778, 30930936, 61997323,
              158727274, 242025902, 226213489, 137672988, 244216783, 49675259, 158168844, 182691070}))
  stage_3_butterfly_27 (
    .x_in(stage_2_per_out[54]),
    .y_in(stage_2_per_out[55]),
    .x_out(stage_3_per_in[54]),
    .y_out(stage_3_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({77981460, 233888407, 199633043, 23405380, 142181410, 169182486, 160841949, 254132077,
              8411857, 34256894, 100229847, 79136411, 75073484, 109479656, 13458851, 205525433,
              192832423, 60548134, 56246211, 140366124, 62117518, 210734246, 148390399, 149992379,
              209085090, 50986641, 10003248, 114486793, 241313184, 266671862, 25944135, 184310992,
              212802310, 237102043, 50222736, 131023241, 18298478, 229100654, 209886001, 196522490,
              145034471, 185138250, 186841927, 122332647, 160807241, 247289727, 258257144, 196328787,
              193915204, 154421517, 92650808, 238382196, 171362072, 171541778, 30930936, 61997323,
              158727274, 242025902, 226213489, 137672988, 244216783, 49675259, 158168844, 182691070}))
  stage_3_butterfly_28 (
    .x_in(stage_2_per_out[56]),
    .y_in(stage_2_per_out[57]),
    .x_out(stage_3_per_in[56]),
    .y_out(stage_3_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({77981460, 233888407, 199633043, 23405380, 142181410, 169182486, 160841949, 254132077,
              8411857, 34256894, 100229847, 79136411, 75073484, 109479656, 13458851, 205525433,
              192832423, 60548134, 56246211, 140366124, 62117518, 210734246, 148390399, 149992379,
              209085090, 50986641, 10003248, 114486793, 241313184, 266671862, 25944135, 184310992,
              212802310, 237102043, 50222736, 131023241, 18298478, 229100654, 209886001, 196522490,
              145034471, 185138250, 186841927, 122332647, 160807241, 247289727, 258257144, 196328787,
              193915204, 154421517, 92650808, 238382196, 171362072, 171541778, 30930936, 61997323,
              158727274, 242025902, 226213489, 137672988, 244216783, 49675259, 158168844, 182691070}))
  stage_3_butterfly_29 (
    .x_in(stage_2_per_out[58]),
    .y_in(stage_2_per_out[59]),
    .x_out(stage_3_per_in[58]),
    .y_out(stage_3_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({77981460, 233888407, 199633043, 23405380, 142181410, 169182486, 160841949, 254132077,
              8411857, 34256894, 100229847, 79136411, 75073484, 109479656, 13458851, 205525433,
              192832423, 60548134, 56246211, 140366124, 62117518, 210734246, 148390399, 149992379,
              209085090, 50986641, 10003248, 114486793, 241313184, 266671862, 25944135, 184310992,
              212802310, 237102043, 50222736, 131023241, 18298478, 229100654, 209886001, 196522490,
              145034471, 185138250, 186841927, 122332647, 160807241, 247289727, 258257144, 196328787,
              193915204, 154421517, 92650808, 238382196, 171362072, 171541778, 30930936, 61997323,
              158727274, 242025902, 226213489, 137672988, 244216783, 49675259, 158168844, 182691070}))
  stage_3_butterfly_30 (
    .x_in(stage_2_per_out[60]),
    .y_in(stage_2_per_out[61]),
    .x_out(stage_3_per_in[60]),
    .y_out(stage_3_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({77981460, 233888407, 199633043, 23405380, 142181410, 169182486, 160841949, 254132077,
              8411857, 34256894, 100229847, 79136411, 75073484, 109479656, 13458851, 205525433,
              192832423, 60548134, 56246211, 140366124, 62117518, 210734246, 148390399, 149992379,
              209085090, 50986641, 10003248, 114486793, 241313184, 266671862, 25944135, 184310992,
              212802310, 237102043, 50222736, 131023241, 18298478, 229100654, 209886001, 196522490,
              145034471, 185138250, 186841927, 122332647, 160807241, 247289727, 258257144, 196328787,
              193915204, 154421517, 92650808, 238382196, 171362072, 171541778, 30930936, 61997323,
              158727274, 242025902, 226213489, 137672988, 244216783, 49675259, 158168844, 182691070}))
  stage_3_butterfly_31 (
    .x_in(stage_2_per_out[62]),
    .y_in(stage_2_per_out[63]),
    .x_out(stage_3_per_in[62]),
    .y_out(stage_3_per_in[63]),
    .clk(clk),
    .rst(rst)
  );




  // TODO(Yang): stage 3 -> stage 4 permutation
  // FIXME: ignore butterfly units for now.
  stage_3_permutation #(
    .DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    .INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_3_4_per (
    .inData_0(stage_3_per_in[0]),
    .inData_1(stage_3_per_in[1]),
    .inData_2(stage_3_per_in[2]),
    .inData_3(stage_3_per_in[3]),
    .inData_4(stage_3_per_in[4]),
    .inData_5(stage_3_per_in[5]),
    .inData_6(stage_3_per_in[6]),
    .inData_7(stage_3_per_in[7]),
    .inData_8(stage_3_per_in[8]),
    .inData_9(stage_3_per_in[9]),
    .inData_10(stage_3_per_in[10]),
    .inData_11(stage_3_per_in[11]),
    .inData_12(stage_3_per_in[12]),
    .inData_13(stage_3_per_in[13]),
    .inData_14(stage_3_per_in[14]),
    .inData_15(stage_3_per_in[15]),
    .inData_16(stage_3_per_in[16]),
    .inData_17(stage_3_per_in[17]),
    .inData_18(stage_3_per_in[18]),
    .inData_19(stage_3_per_in[19]),
    .inData_20(stage_3_per_in[20]),
    .inData_21(stage_3_per_in[21]),
    .inData_22(stage_3_per_in[22]),
    .inData_23(stage_3_per_in[23]),
    .inData_24(stage_3_per_in[24]),
    .inData_25(stage_3_per_in[25]),
    .inData_26(stage_3_per_in[26]),
    .inData_27(stage_3_per_in[27]),
    .inData_28(stage_3_per_in[28]),
    .inData_29(stage_3_per_in[29]),
    .inData_30(stage_3_per_in[30]),
    .inData_31(stage_3_per_in[31]),
    .inData_32(stage_3_per_in[32]),
    .inData_33(stage_3_per_in[33]),
    .inData_34(stage_3_per_in[34]),
    .inData_35(stage_3_per_in[35]),
    .inData_36(stage_3_per_in[36]),
    .inData_37(stage_3_per_in[37]),
    .inData_38(stage_3_per_in[38]),
    .inData_39(stage_3_per_in[39]),
    .inData_40(stage_3_per_in[40]),
    .inData_41(stage_3_per_in[41]),
    .inData_42(stage_3_per_in[42]),
    .inData_43(stage_3_per_in[43]),
    .inData_44(stage_3_per_in[44]),
    .inData_45(stage_3_per_in[45]),
    .inData_46(stage_3_per_in[46]),
    .inData_47(stage_3_per_in[47]),
    .inData_48(stage_3_per_in[48]),
    .inData_49(stage_3_per_in[49]),
    .inData_50(stage_3_per_in[50]),
    .inData_51(stage_3_per_in[51]),
    .inData_52(stage_3_per_in[52]),
    .inData_53(stage_3_per_in[53]),
    .inData_54(stage_3_per_in[54]),
    .inData_55(stage_3_per_in[55]),
    .inData_56(stage_3_per_in[56]),
    .inData_57(stage_3_per_in[57]),
    .inData_58(stage_3_per_in[58]),
    .inData_59(stage_3_per_in[59]),
    .inData_60(stage_3_per_in[60]),
    .inData_61(stage_3_per_in[61]),
    .inData_62(stage_3_per_in[62]),
    .inData_63(stage_3_per_in[63]),
    .outData_0(stage_3_per_out[0]),
    .outData_1(stage_3_per_out[1]),
    .outData_2(stage_3_per_out[2]),
    .outData_3(stage_3_per_out[3]),
    .outData_4(stage_3_per_out[4]),
    .outData_5(stage_3_per_out[5]),
    .outData_6(stage_3_per_out[6]),
    .outData_7(stage_3_per_out[7]),
    .outData_8(stage_3_per_out[8]),
    .outData_9(stage_3_per_out[9]),
    .outData_10(stage_3_per_out[10]),
    .outData_11(stage_3_per_out[11]),
    .outData_12(stage_3_per_out[12]),
    .outData_13(stage_3_per_out[13]),
    .outData_14(stage_3_per_out[14]),
    .outData_15(stage_3_per_out[15]),
    .outData_16(stage_3_per_out[16]),
    .outData_17(stage_3_per_out[17]),
    .outData_18(stage_3_per_out[18]),
    .outData_19(stage_3_per_out[19]),
    .outData_20(stage_3_per_out[20]),
    .outData_21(stage_3_per_out[21]),
    .outData_22(stage_3_per_out[22]),
    .outData_23(stage_3_per_out[23]),
    .outData_24(stage_3_per_out[24]),
    .outData_25(stage_3_per_out[25]),
    .outData_26(stage_3_per_out[26]),
    .outData_27(stage_3_per_out[27]),
    .outData_28(stage_3_per_out[28]),
    .outData_29(stage_3_per_out[29]),
    .outData_30(stage_3_per_out[30]),
    .outData_31(stage_3_per_out[31]),
    .outData_32(stage_3_per_out[32]),
    .outData_33(stage_3_per_out[33]),
    .outData_34(stage_3_per_out[34]),
    .outData_35(stage_3_per_out[35]),
    .outData_36(stage_3_per_out[36]),
    .outData_37(stage_3_per_out[37]),
    .outData_38(stage_3_per_out[38]),
    .outData_39(stage_3_per_out[39]),
    .outData_40(stage_3_per_out[40]),
    .outData_41(stage_3_per_out[41]),
    .outData_42(stage_3_per_out[42]),
    .outData_43(stage_3_per_out[43]),
    .outData_44(stage_3_per_out[44]),
    .outData_45(stage_3_per_out[45]),
    .outData_46(stage_3_per_out[46]),
    .outData_47(stage_3_per_out[47]),
    .outData_48(stage_3_per_out[48]),
    .outData_49(stage_3_per_out[49]),
    .outData_50(stage_3_per_out[50]),
    .outData_51(stage_3_per_out[51]),
    .outData_52(stage_3_per_out[52]),
    .outData_53(stage_3_per_out[53]),
    .outData_54(stage_3_per_out[54]),
    .outData_55(stage_3_per_out[55]),
    .outData_56(stage_3_per_out[56]),
    .outData_57(stage_3_per_out[57]),
    .outData_58(stage_3_per_out[58]),
    .outData_59(stage_3_per_out[59]),
    .outData_60(stage_3_per_out[60]),
    .outData_61(stage_3_per_out[61]),
    .outData_62(stage_3_per_out[62]),
    .outData_63(stage_3_per_out[63]),
    .in_start(in_start[3]),
    .out_start(out_start[3]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 4 32 butterfly units
  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 116401819, 11101448, 71064168, 189762285, 81956368, 244883276, 135288005,
              229228230, 216143425, 101839787, 265950570, 85922744, 254450415, 10571783, 14542514,
              117496916, 250166212, 192696288, 130557622, 106640438, 234030247, 90597117, 209086118,
              189881206, 10130658, 241125460, 176471684, 209161759, 231358848, 245906264, 63350037,
              55721255, 47751177, 64217206, 229216409, 40553702, 204666342, 214551729, 33479018,
              226739459, 34119889, 246744565, 2795054, 104557084, 96142103, 104784816, 41086336,
              122008382, 211668928, 225636920, 197074908, 47994339, 252442032, 168407516, 9720223,
              184226747, 143969713, 69161747, 245828202, 239545014, 98878775, 72738487, 217644581}))
  stage_4_butterfly_0 (
    .x_in(stage_3_per_out[0]),
    .y_in(stage_3_per_out[1]),
    .x_out(stage_4_per_in[0]),
    .y_out(stage_4_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 116401819, 11101448, 71064168, 189762285, 81956368, 244883276, 135288005,
              229228230, 216143425, 101839787, 265950570, 85922744, 254450415, 10571783, 14542514,
              117496916, 250166212, 192696288, 130557622, 106640438, 234030247, 90597117, 209086118,
              189881206, 10130658, 241125460, 176471684, 209161759, 231358848, 245906264, 63350037,
              55721255, 47751177, 64217206, 229216409, 40553702, 204666342, 214551729, 33479018,
              226739459, 34119889, 246744565, 2795054, 104557084, 96142103, 104784816, 41086336,
              122008382, 211668928, 225636920, 197074908, 47994339, 252442032, 168407516, 9720223,
              184226747, 143969713, 69161747, 245828202, 239545014, 98878775, 72738487, 217644581}))
  stage_4_butterfly_1 (
    .x_in(stage_3_per_out[2]),
    .y_in(stage_3_per_out[3]),
    .x_out(stage_4_per_in[2]),
    .y_out(stage_4_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 116401819, 11101448, 71064168, 189762285, 81956368, 244883276, 135288005,
              229228230, 216143425, 101839787, 265950570, 85922744, 254450415, 10571783, 14542514,
              117496916, 250166212, 192696288, 130557622, 106640438, 234030247, 90597117, 209086118,
              189881206, 10130658, 241125460, 176471684, 209161759, 231358848, 245906264, 63350037,
              55721255, 47751177, 64217206, 229216409, 40553702, 204666342, 214551729, 33479018,
              226739459, 34119889, 246744565, 2795054, 104557084, 96142103, 104784816, 41086336,
              122008382, 211668928, 225636920, 197074908, 47994339, 252442032, 168407516, 9720223,
              184226747, 143969713, 69161747, 245828202, 239545014, 98878775, 72738487, 217644581}))
  stage_4_butterfly_2 (
    .x_in(stage_3_per_out[4]),
    .y_in(stage_3_per_out[5]),
    .x_out(stage_4_per_in[4]),
    .y_out(stage_4_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 116401819, 11101448, 71064168, 189762285, 81956368, 244883276, 135288005,
              229228230, 216143425, 101839787, 265950570, 85922744, 254450415, 10571783, 14542514,
              117496916, 250166212, 192696288, 130557622, 106640438, 234030247, 90597117, 209086118,
              189881206, 10130658, 241125460, 176471684, 209161759, 231358848, 245906264, 63350037,
              55721255, 47751177, 64217206, 229216409, 40553702, 204666342, 214551729, 33479018,
              226739459, 34119889, 246744565, 2795054, 104557084, 96142103, 104784816, 41086336,
              122008382, 211668928, 225636920, 197074908, 47994339, 252442032, 168407516, 9720223,
              184226747, 143969713, 69161747, 245828202, 239545014, 98878775, 72738487, 217644581}))
  stage_4_butterfly_3 (
    .x_in(stage_3_per_out[6]),
    .y_in(stage_3_per_out[7]),
    .x_out(stage_4_per_in[6]),
    .y_out(stage_4_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 116401819, 11101448, 71064168, 189762285, 81956368, 244883276, 135288005,
              229228230, 216143425, 101839787, 265950570, 85922744, 254450415, 10571783, 14542514,
              117496916, 250166212, 192696288, 130557622, 106640438, 234030247, 90597117, 209086118,
              189881206, 10130658, 241125460, 176471684, 209161759, 231358848, 245906264, 63350037,
              55721255, 47751177, 64217206, 229216409, 40553702, 204666342, 214551729, 33479018,
              226739459, 34119889, 246744565, 2795054, 104557084, 96142103, 104784816, 41086336,
              122008382, 211668928, 225636920, 197074908, 47994339, 252442032, 168407516, 9720223,
              184226747, 143969713, 69161747, 245828202, 239545014, 98878775, 72738487, 217644581}))
  stage_4_butterfly_4 (
    .x_in(stage_3_per_out[8]),
    .y_in(stage_3_per_out[9]),
    .x_out(stage_4_per_in[8]),
    .y_out(stage_4_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 116401819, 11101448, 71064168, 189762285, 81956368, 244883276, 135288005,
              229228230, 216143425, 101839787, 265950570, 85922744, 254450415, 10571783, 14542514,
              117496916, 250166212, 192696288, 130557622, 106640438, 234030247, 90597117, 209086118,
              189881206, 10130658, 241125460, 176471684, 209161759, 231358848, 245906264, 63350037,
              55721255, 47751177, 64217206, 229216409, 40553702, 204666342, 214551729, 33479018,
              226739459, 34119889, 246744565, 2795054, 104557084, 96142103, 104784816, 41086336,
              122008382, 211668928, 225636920, 197074908, 47994339, 252442032, 168407516, 9720223,
              184226747, 143969713, 69161747, 245828202, 239545014, 98878775, 72738487, 217644581}))
  stage_4_butterfly_5 (
    .x_in(stage_3_per_out[10]),
    .y_in(stage_3_per_out[11]),
    .x_out(stage_4_per_in[10]),
    .y_out(stage_4_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 116401819, 11101448, 71064168, 189762285, 81956368, 244883276, 135288005,
              229228230, 216143425, 101839787, 265950570, 85922744, 254450415, 10571783, 14542514,
              117496916, 250166212, 192696288, 130557622, 106640438, 234030247, 90597117, 209086118,
              189881206, 10130658, 241125460, 176471684, 209161759, 231358848, 245906264, 63350037,
              55721255, 47751177, 64217206, 229216409, 40553702, 204666342, 214551729, 33479018,
              226739459, 34119889, 246744565, 2795054, 104557084, 96142103, 104784816, 41086336,
              122008382, 211668928, 225636920, 197074908, 47994339, 252442032, 168407516, 9720223,
              184226747, 143969713, 69161747, 245828202, 239545014, 98878775, 72738487, 217644581}))
  stage_4_butterfly_6 (
    .x_in(stage_3_per_out[12]),
    .y_in(stage_3_per_out[13]),
    .x_out(stage_4_per_in[12]),
    .y_out(stage_4_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 116401819, 11101448, 71064168, 189762285, 81956368, 244883276, 135288005,
              229228230, 216143425, 101839787, 265950570, 85922744, 254450415, 10571783, 14542514,
              117496916, 250166212, 192696288, 130557622, 106640438, 234030247, 90597117, 209086118,
              189881206, 10130658, 241125460, 176471684, 209161759, 231358848, 245906264, 63350037,
              55721255, 47751177, 64217206, 229216409, 40553702, 204666342, 214551729, 33479018,
              226739459, 34119889, 246744565, 2795054, 104557084, 96142103, 104784816, 41086336,
              122008382, 211668928, 225636920, 197074908, 47994339, 252442032, 168407516, 9720223,
              184226747, 143969713, 69161747, 245828202, 239545014, 98878775, 72738487, 217644581}))
  stage_4_butterfly_7 (
    .x_in(stage_3_per_out[14]),
    .y_in(stage_3_per_out[15]),
    .x_out(stage_4_per_in[14]),
    .y_out(stage_4_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 116401819, 11101448, 71064168, 189762285, 81956368, 244883276, 135288005,
              229228230, 216143425, 101839787, 265950570, 85922744, 254450415, 10571783, 14542514,
              117496916, 250166212, 192696288, 130557622, 106640438, 234030247, 90597117, 209086118,
              189881206, 10130658, 241125460, 176471684, 209161759, 231358848, 245906264, 63350037,
              55721255, 47751177, 64217206, 229216409, 40553702, 204666342, 214551729, 33479018,
              226739459, 34119889, 246744565, 2795054, 104557084, 96142103, 104784816, 41086336,
              122008382, 211668928, 225636920, 197074908, 47994339, 252442032, 168407516, 9720223,
              184226747, 143969713, 69161747, 245828202, 239545014, 98878775, 72738487, 217644581}))
  stage_4_butterfly_8 (
    .x_in(stage_3_per_out[16]),
    .y_in(stage_3_per_out[17]),
    .x_out(stage_4_per_in[16]),
    .y_out(stage_4_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 116401819, 11101448, 71064168, 189762285, 81956368, 244883276, 135288005,
              229228230, 216143425, 101839787, 265950570, 85922744, 254450415, 10571783, 14542514,
              117496916, 250166212, 192696288, 130557622, 106640438, 234030247, 90597117, 209086118,
              189881206, 10130658, 241125460, 176471684, 209161759, 231358848, 245906264, 63350037,
              55721255, 47751177, 64217206, 229216409, 40553702, 204666342, 214551729, 33479018,
              226739459, 34119889, 246744565, 2795054, 104557084, 96142103, 104784816, 41086336,
              122008382, 211668928, 225636920, 197074908, 47994339, 252442032, 168407516, 9720223,
              184226747, 143969713, 69161747, 245828202, 239545014, 98878775, 72738487, 217644581}))
  stage_4_butterfly_9 (
    .x_in(stage_3_per_out[18]),
    .y_in(stage_3_per_out[19]),
    .x_out(stage_4_per_in[18]),
    .y_out(stage_4_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 116401819, 11101448, 71064168, 189762285, 81956368, 244883276, 135288005,
              229228230, 216143425, 101839787, 265950570, 85922744, 254450415, 10571783, 14542514,
              117496916, 250166212, 192696288, 130557622, 106640438, 234030247, 90597117, 209086118,
              189881206, 10130658, 241125460, 176471684, 209161759, 231358848, 245906264, 63350037,
              55721255, 47751177, 64217206, 229216409, 40553702, 204666342, 214551729, 33479018,
              226739459, 34119889, 246744565, 2795054, 104557084, 96142103, 104784816, 41086336,
              122008382, 211668928, 225636920, 197074908, 47994339, 252442032, 168407516, 9720223,
              184226747, 143969713, 69161747, 245828202, 239545014, 98878775, 72738487, 217644581}))
  stage_4_butterfly_10 (
    .x_in(stage_3_per_out[20]),
    .y_in(stage_3_per_out[21]),
    .x_out(stage_4_per_in[20]),
    .y_out(stage_4_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 116401819, 11101448, 71064168, 189762285, 81956368, 244883276, 135288005,
              229228230, 216143425, 101839787, 265950570, 85922744, 254450415, 10571783, 14542514,
              117496916, 250166212, 192696288, 130557622, 106640438, 234030247, 90597117, 209086118,
              189881206, 10130658, 241125460, 176471684, 209161759, 231358848, 245906264, 63350037,
              55721255, 47751177, 64217206, 229216409, 40553702, 204666342, 214551729, 33479018,
              226739459, 34119889, 246744565, 2795054, 104557084, 96142103, 104784816, 41086336,
              122008382, 211668928, 225636920, 197074908, 47994339, 252442032, 168407516, 9720223,
              184226747, 143969713, 69161747, 245828202, 239545014, 98878775, 72738487, 217644581}))
  stage_4_butterfly_11 (
    .x_in(stage_3_per_out[22]),
    .y_in(stage_3_per_out[23]),
    .x_out(stage_4_per_in[22]),
    .y_out(stage_4_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 116401819, 11101448, 71064168, 189762285, 81956368, 244883276, 135288005,
              229228230, 216143425, 101839787, 265950570, 85922744, 254450415, 10571783, 14542514,
              117496916, 250166212, 192696288, 130557622, 106640438, 234030247, 90597117, 209086118,
              189881206, 10130658, 241125460, 176471684, 209161759, 231358848, 245906264, 63350037,
              55721255, 47751177, 64217206, 229216409, 40553702, 204666342, 214551729, 33479018,
              226739459, 34119889, 246744565, 2795054, 104557084, 96142103, 104784816, 41086336,
              122008382, 211668928, 225636920, 197074908, 47994339, 252442032, 168407516, 9720223,
              184226747, 143969713, 69161747, 245828202, 239545014, 98878775, 72738487, 217644581}))
  stage_4_butterfly_12 (
    .x_in(stage_3_per_out[24]),
    .y_in(stage_3_per_out[25]),
    .x_out(stage_4_per_in[24]),
    .y_out(stage_4_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 116401819, 11101448, 71064168, 189762285, 81956368, 244883276, 135288005,
              229228230, 216143425, 101839787, 265950570, 85922744, 254450415, 10571783, 14542514,
              117496916, 250166212, 192696288, 130557622, 106640438, 234030247, 90597117, 209086118,
              189881206, 10130658, 241125460, 176471684, 209161759, 231358848, 245906264, 63350037,
              55721255, 47751177, 64217206, 229216409, 40553702, 204666342, 214551729, 33479018,
              226739459, 34119889, 246744565, 2795054, 104557084, 96142103, 104784816, 41086336,
              122008382, 211668928, 225636920, 197074908, 47994339, 252442032, 168407516, 9720223,
              184226747, 143969713, 69161747, 245828202, 239545014, 98878775, 72738487, 217644581}))
  stage_4_butterfly_13 (
    .x_in(stage_3_per_out[26]),
    .y_in(stage_3_per_out[27]),
    .x_out(stage_4_per_in[26]),
    .y_out(stage_4_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 116401819, 11101448, 71064168, 189762285, 81956368, 244883276, 135288005,
              229228230, 216143425, 101839787, 265950570, 85922744, 254450415, 10571783, 14542514,
              117496916, 250166212, 192696288, 130557622, 106640438, 234030247, 90597117, 209086118,
              189881206, 10130658, 241125460, 176471684, 209161759, 231358848, 245906264, 63350037,
              55721255, 47751177, 64217206, 229216409, 40553702, 204666342, 214551729, 33479018,
              226739459, 34119889, 246744565, 2795054, 104557084, 96142103, 104784816, 41086336,
              122008382, 211668928, 225636920, 197074908, 47994339, 252442032, 168407516, 9720223,
              184226747, 143969713, 69161747, 245828202, 239545014, 98878775, 72738487, 217644581}))
  stage_4_butterfly_14 (
    .x_in(stage_3_per_out[28]),
    .y_in(stage_3_per_out[29]),
    .x_out(stage_4_per_in[28]),
    .y_out(stage_4_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 116401819, 11101448, 71064168, 189762285, 81956368, 244883276, 135288005,
              229228230, 216143425, 101839787, 265950570, 85922744, 254450415, 10571783, 14542514,
              117496916, 250166212, 192696288, 130557622, 106640438, 234030247, 90597117, 209086118,
              189881206, 10130658, 241125460, 176471684, 209161759, 231358848, 245906264, 63350037,
              55721255, 47751177, 64217206, 229216409, 40553702, 204666342, 214551729, 33479018,
              226739459, 34119889, 246744565, 2795054, 104557084, 96142103, 104784816, 41086336,
              122008382, 211668928, 225636920, 197074908, 47994339, 252442032, 168407516, 9720223,
              184226747, 143969713, 69161747, 245828202, 239545014, 98878775, 72738487, 217644581}))
  stage_4_butterfly_15 (
    .x_in(stage_3_per_out[30]),
    .y_in(stage_3_per_out[31]),
    .x_out(stage_4_per_in[30]),
    .y_out(stage_4_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 18729522, 68136911, 166886297, 21713495, 176917280, 7055647, 238498066,
              148662095, 181639510, 256040960, 240677074, 123185272, 97765534, 170227406, 40475021,
              193371292, 167885779, 159404461, 37051834, 183348420, 41155851, 173702965, 258612781,
              186592442, 139182289, 243304319, 83853696, 236144340, 230433664, 189591954, 54284329,
              254509489, 15417588, 66148505, 108083129, 118518376, 241682233, 108810259, 223427563,
              67012048, 77337691, 104174682, 161827885, 155168409, 118841873, 3883583, 134866823,
              25569479, 123954975, 120936039, 210298252, 13519489, 162031725, 132703565, 19493867,
              71933862, 230702770, 180525688, 13250338, 139555205, 9446767, 171721518, 249970613}))
  stage_4_butterfly_16 (
    .x_in(stage_3_per_out[32]),
    .y_in(stage_3_per_out[33]),
    .x_out(stage_4_per_in[32]),
    .y_out(stage_4_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 18729522, 68136911, 166886297, 21713495, 176917280, 7055647, 238498066,
              148662095, 181639510, 256040960, 240677074, 123185272, 97765534, 170227406, 40475021,
              193371292, 167885779, 159404461, 37051834, 183348420, 41155851, 173702965, 258612781,
              186592442, 139182289, 243304319, 83853696, 236144340, 230433664, 189591954, 54284329,
              254509489, 15417588, 66148505, 108083129, 118518376, 241682233, 108810259, 223427563,
              67012048, 77337691, 104174682, 161827885, 155168409, 118841873, 3883583, 134866823,
              25569479, 123954975, 120936039, 210298252, 13519489, 162031725, 132703565, 19493867,
              71933862, 230702770, 180525688, 13250338, 139555205, 9446767, 171721518, 249970613}))
  stage_4_butterfly_17 (
    .x_in(stage_3_per_out[34]),
    .y_in(stage_3_per_out[35]),
    .x_out(stage_4_per_in[34]),
    .y_out(stage_4_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 18729522, 68136911, 166886297, 21713495, 176917280, 7055647, 238498066,
              148662095, 181639510, 256040960, 240677074, 123185272, 97765534, 170227406, 40475021,
              193371292, 167885779, 159404461, 37051834, 183348420, 41155851, 173702965, 258612781,
              186592442, 139182289, 243304319, 83853696, 236144340, 230433664, 189591954, 54284329,
              254509489, 15417588, 66148505, 108083129, 118518376, 241682233, 108810259, 223427563,
              67012048, 77337691, 104174682, 161827885, 155168409, 118841873, 3883583, 134866823,
              25569479, 123954975, 120936039, 210298252, 13519489, 162031725, 132703565, 19493867,
              71933862, 230702770, 180525688, 13250338, 139555205, 9446767, 171721518, 249970613}))
  stage_4_butterfly_18 (
    .x_in(stage_3_per_out[36]),
    .y_in(stage_3_per_out[37]),
    .x_out(stage_4_per_in[36]),
    .y_out(stage_4_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 18729522, 68136911, 166886297, 21713495, 176917280, 7055647, 238498066,
              148662095, 181639510, 256040960, 240677074, 123185272, 97765534, 170227406, 40475021,
              193371292, 167885779, 159404461, 37051834, 183348420, 41155851, 173702965, 258612781,
              186592442, 139182289, 243304319, 83853696, 236144340, 230433664, 189591954, 54284329,
              254509489, 15417588, 66148505, 108083129, 118518376, 241682233, 108810259, 223427563,
              67012048, 77337691, 104174682, 161827885, 155168409, 118841873, 3883583, 134866823,
              25569479, 123954975, 120936039, 210298252, 13519489, 162031725, 132703565, 19493867,
              71933862, 230702770, 180525688, 13250338, 139555205, 9446767, 171721518, 249970613}))
  stage_4_butterfly_19 (
    .x_in(stage_3_per_out[38]),
    .y_in(stage_3_per_out[39]),
    .x_out(stage_4_per_in[38]),
    .y_out(stage_4_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 18729522, 68136911, 166886297, 21713495, 176917280, 7055647, 238498066,
              148662095, 181639510, 256040960, 240677074, 123185272, 97765534, 170227406, 40475021,
              193371292, 167885779, 159404461, 37051834, 183348420, 41155851, 173702965, 258612781,
              186592442, 139182289, 243304319, 83853696, 236144340, 230433664, 189591954, 54284329,
              254509489, 15417588, 66148505, 108083129, 118518376, 241682233, 108810259, 223427563,
              67012048, 77337691, 104174682, 161827885, 155168409, 118841873, 3883583, 134866823,
              25569479, 123954975, 120936039, 210298252, 13519489, 162031725, 132703565, 19493867,
              71933862, 230702770, 180525688, 13250338, 139555205, 9446767, 171721518, 249970613}))
  stage_4_butterfly_20 (
    .x_in(stage_3_per_out[40]),
    .y_in(stage_3_per_out[41]),
    .x_out(stage_4_per_in[40]),
    .y_out(stage_4_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 18729522, 68136911, 166886297, 21713495, 176917280, 7055647, 238498066,
              148662095, 181639510, 256040960, 240677074, 123185272, 97765534, 170227406, 40475021,
              193371292, 167885779, 159404461, 37051834, 183348420, 41155851, 173702965, 258612781,
              186592442, 139182289, 243304319, 83853696, 236144340, 230433664, 189591954, 54284329,
              254509489, 15417588, 66148505, 108083129, 118518376, 241682233, 108810259, 223427563,
              67012048, 77337691, 104174682, 161827885, 155168409, 118841873, 3883583, 134866823,
              25569479, 123954975, 120936039, 210298252, 13519489, 162031725, 132703565, 19493867,
              71933862, 230702770, 180525688, 13250338, 139555205, 9446767, 171721518, 249970613}))
  stage_4_butterfly_21 (
    .x_in(stage_3_per_out[42]),
    .y_in(stage_3_per_out[43]),
    .x_out(stage_4_per_in[42]),
    .y_out(stage_4_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 18729522, 68136911, 166886297, 21713495, 176917280, 7055647, 238498066,
              148662095, 181639510, 256040960, 240677074, 123185272, 97765534, 170227406, 40475021,
              193371292, 167885779, 159404461, 37051834, 183348420, 41155851, 173702965, 258612781,
              186592442, 139182289, 243304319, 83853696, 236144340, 230433664, 189591954, 54284329,
              254509489, 15417588, 66148505, 108083129, 118518376, 241682233, 108810259, 223427563,
              67012048, 77337691, 104174682, 161827885, 155168409, 118841873, 3883583, 134866823,
              25569479, 123954975, 120936039, 210298252, 13519489, 162031725, 132703565, 19493867,
              71933862, 230702770, 180525688, 13250338, 139555205, 9446767, 171721518, 249970613}))
  stage_4_butterfly_22 (
    .x_in(stage_3_per_out[44]),
    .y_in(stage_3_per_out[45]),
    .x_out(stage_4_per_in[44]),
    .y_out(stage_4_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 18729522, 68136911, 166886297, 21713495, 176917280, 7055647, 238498066,
              148662095, 181639510, 256040960, 240677074, 123185272, 97765534, 170227406, 40475021,
              193371292, 167885779, 159404461, 37051834, 183348420, 41155851, 173702965, 258612781,
              186592442, 139182289, 243304319, 83853696, 236144340, 230433664, 189591954, 54284329,
              254509489, 15417588, 66148505, 108083129, 118518376, 241682233, 108810259, 223427563,
              67012048, 77337691, 104174682, 161827885, 155168409, 118841873, 3883583, 134866823,
              25569479, 123954975, 120936039, 210298252, 13519489, 162031725, 132703565, 19493867,
              71933862, 230702770, 180525688, 13250338, 139555205, 9446767, 171721518, 249970613}))
  stage_4_butterfly_23 (
    .x_in(stage_3_per_out[46]),
    .y_in(stage_3_per_out[47]),
    .x_out(stage_4_per_in[46]),
    .y_out(stage_4_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 18729522, 68136911, 166886297, 21713495, 176917280, 7055647, 238498066,
              148662095, 181639510, 256040960, 240677074, 123185272, 97765534, 170227406, 40475021,
              193371292, 167885779, 159404461, 37051834, 183348420, 41155851, 173702965, 258612781,
              186592442, 139182289, 243304319, 83853696, 236144340, 230433664, 189591954, 54284329,
              254509489, 15417588, 66148505, 108083129, 118518376, 241682233, 108810259, 223427563,
              67012048, 77337691, 104174682, 161827885, 155168409, 118841873, 3883583, 134866823,
              25569479, 123954975, 120936039, 210298252, 13519489, 162031725, 132703565, 19493867,
              71933862, 230702770, 180525688, 13250338, 139555205, 9446767, 171721518, 249970613}))
  stage_4_butterfly_24 (
    .x_in(stage_3_per_out[48]),
    .y_in(stage_3_per_out[49]),
    .x_out(stage_4_per_in[48]),
    .y_out(stage_4_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 18729522, 68136911, 166886297, 21713495, 176917280, 7055647, 238498066,
              148662095, 181639510, 256040960, 240677074, 123185272, 97765534, 170227406, 40475021,
              193371292, 167885779, 159404461, 37051834, 183348420, 41155851, 173702965, 258612781,
              186592442, 139182289, 243304319, 83853696, 236144340, 230433664, 189591954, 54284329,
              254509489, 15417588, 66148505, 108083129, 118518376, 241682233, 108810259, 223427563,
              67012048, 77337691, 104174682, 161827885, 155168409, 118841873, 3883583, 134866823,
              25569479, 123954975, 120936039, 210298252, 13519489, 162031725, 132703565, 19493867,
              71933862, 230702770, 180525688, 13250338, 139555205, 9446767, 171721518, 249970613}))
  stage_4_butterfly_25 (
    .x_in(stage_3_per_out[50]),
    .y_in(stage_3_per_out[51]),
    .x_out(stage_4_per_in[50]),
    .y_out(stage_4_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 18729522, 68136911, 166886297, 21713495, 176917280, 7055647, 238498066,
              148662095, 181639510, 256040960, 240677074, 123185272, 97765534, 170227406, 40475021,
              193371292, 167885779, 159404461, 37051834, 183348420, 41155851, 173702965, 258612781,
              186592442, 139182289, 243304319, 83853696, 236144340, 230433664, 189591954, 54284329,
              254509489, 15417588, 66148505, 108083129, 118518376, 241682233, 108810259, 223427563,
              67012048, 77337691, 104174682, 161827885, 155168409, 118841873, 3883583, 134866823,
              25569479, 123954975, 120936039, 210298252, 13519489, 162031725, 132703565, 19493867,
              71933862, 230702770, 180525688, 13250338, 139555205, 9446767, 171721518, 249970613}))
  stage_4_butterfly_26 (
    .x_in(stage_3_per_out[52]),
    .y_in(stage_3_per_out[53]),
    .x_out(stage_4_per_in[52]),
    .y_out(stage_4_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 18729522, 68136911, 166886297, 21713495, 176917280, 7055647, 238498066,
              148662095, 181639510, 256040960, 240677074, 123185272, 97765534, 170227406, 40475021,
              193371292, 167885779, 159404461, 37051834, 183348420, 41155851, 173702965, 258612781,
              186592442, 139182289, 243304319, 83853696, 236144340, 230433664, 189591954, 54284329,
              254509489, 15417588, 66148505, 108083129, 118518376, 241682233, 108810259, 223427563,
              67012048, 77337691, 104174682, 161827885, 155168409, 118841873, 3883583, 134866823,
              25569479, 123954975, 120936039, 210298252, 13519489, 162031725, 132703565, 19493867,
              71933862, 230702770, 180525688, 13250338, 139555205, 9446767, 171721518, 249970613}))
  stage_4_butterfly_27 (
    .x_in(stage_3_per_out[54]),
    .y_in(stage_3_per_out[55]),
    .x_out(stage_4_per_in[54]),
    .y_out(stage_4_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 18729522, 68136911, 166886297, 21713495, 176917280, 7055647, 238498066,
              148662095, 181639510, 256040960, 240677074, 123185272, 97765534, 170227406, 40475021,
              193371292, 167885779, 159404461, 37051834, 183348420, 41155851, 173702965, 258612781,
              186592442, 139182289, 243304319, 83853696, 236144340, 230433664, 189591954, 54284329,
              254509489, 15417588, 66148505, 108083129, 118518376, 241682233, 108810259, 223427563,
              67012048, 77337691, 104174682, 161827885, 155168409, 118841873, 3883583, 134866823,
              25569479, 123954975, 120936039, 210298252, 13519489, 162031725, 132703565, 19493867,
              71933862, 230702770, 180525688, 13250338, 139555205, 9446767, 171721518, 249970613}))
  stage_4_butterfly_28 (
    .x_in(stage_3_per_out[56]),
    .y_in(stage_3_per_out[57]),
    .x_out(stage_4_per_in[56]),
    .y_out(stage_4_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 18729522, 68136911, 166886297, 21713495, 176917280, 7055647, 238498066,
              148662095, 181639510, 256040960, 240677074, 123185272, 97765534, 170227406, 40475021,
              193371292, 167885779, 159404461, 37051834, 183348420, 41155851, 173702965, 258612781,
              186592442, 139182289, 243304319, 83853696, 236144340, 230433664, 189591954, 54284329,
              254509489, 15417588, 66148505, 108083129, 118518376, 241682233, 108810259, 223427563,
              67012048, 77337691, 104174682, 161827885, 155168409, 118841873, 3883583, 134866823,
              25569479, 123954975, 120936039, 210298252, 13519489, 162031725, 132703565, 19493867,
              71933862, 230702770, 180525688, 13250338, 139555205, 9446767, 171721518, 249970613}))
  stage_4_butterfly_29 (
    .x_in(stage_3_per_out[58]),
    .y_in(stage_3_per_out[59]),
    .x_out(stage_4_per_in[58]),
    .y_out(stage_4_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 18729522, 68136911, 166886297, 21713495, 176917280, 7055647, 238498066,
              148662095, 181639510, 256040960, 240677074, 123185272, 97765534, 170227406, 40475021,
              193371292, 167885779, 159404461, 37051834, 183348420, 41155851, 173702965, 258612781,
              186592442, 139182289, 243304319, 83853696, 236144340, 230433664, 189591954, 54284329,
              254509489, 15417588, 66148505, 108083129, 118518376, 241682233, 108810259, 223427563,
              67012048, 77337691, 104174682, 161827885, 155168409, 118841873, 3883583, 134866823,
              25569479, 123954975, 120936039, 210298252, 13519489, 162031725, 132703565, 19493867,
              71933862, 230702770, 180525688, 13250338, 139555205, 9446767, 171721518, 249970613}))
  stage_4_butterfly_30 (
    .x_in(stage_3_per_out[60]),
    .y_in(stage_3_per_out[61]),
    .x_out(stage_4_per_in[60]),
    .y_out(stage_4_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 18729522, 68136911, 166886297, 21713495, 176917280, 7055647, 238498066,
              148662095, 181639510, 256040960, 240677074, 123185272, 97765534, 170227406, 40475021,
              193371292, 167885779, 159404461, 37051834, 183348420, 41155851, 173702965, 258612781,
              186592442, 139182289, 243304319, 83853696, 236144340, 230433664, 189591954, 54284329,
              254509489, 15417588, 66148505, 108083129, 118518376, 241682233, 108810259, 223427563,
              67012048, 77337691, 104174682, 161827885, 155168409, 118841873, 3883583, 134866823,
              25569479, 123954975, 120936039, 210298252, 13519489, 162031725, 132703565, 19493867,
              71933862, 230702770, 180525688, 13250338, 139555205, 9446767, 171721518, 249970613}))
  stage_4_butterfly_31 (
    .x_in(stage_3_per_out[62]),
    .y_in(stage_3_per_out[63]),
    .x_out(stage_4_per_in[62]),
    .y_out(stage_4_per_in[63]),
    .clk(clk),
    .rst(rst)
  );



  // TODO(Yang): stage 4 -> stage 5 permutation
  // FIXME: ignore butterfly units for now.
  stage_4_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_4_5_per (
    .inData_0(stage_4_per_in[0]),
    .inData_1(stage_4_per_in[1]),
    .inData_2(stage_4_per_in[2]),
    .inData_3(stage_4_per_in[3]),
    .inData_4(stage_4_per_in[4]),
    .inData_5(stage_4_per_in[5]),
    .inData_6(stage_4_per_in[6]),
    .inData_7(stage_4_per_in[7]),
    .inData_8(stage_4_per_in[8]),
    .inData_9(stage_4_per_in[9]),
    .inData_10(stage_4_per_in[10]),
    .inData_11(stage_4_per_in[11]),
    .inData_12(stage_4_per_in[12]),
    .inData_13(stage_4_per_in[13]),
    .inData_14(stage_4_per_in[14]),
    .inData_15(stage_4_per_in[15]),
    .inData_16(stage_4_per_in[16]),
    .inData_17(stage_4_per_in[17]),
    .inData_18(stage_4_per_in[18]),
    .inData_19(stage_4_per_in[19]),
    .inData_20(stage_4_per_in[20]),
    .inData_21(stage_4_per_in[21]),
    .inData_22(stage_4_per_in[22]),
    .inData_23(stage_4_per_in[23]),
    .inData_24(stage_4_per_in[24]),
    .inData_25(stage_4_per_in[25]),
    .inData_26(stage_4_per_in[26]),
    .inData_27(stage_4_per_in[27]),
    .inData_28(stage_4_per_in[28]),
    .inData_29(stage_4_per_in[29]),
    .inData_30(stage_4_per_in[30]),
    .inData_31(stage_4_per_in[31]),
    .inData_32(stage_4_per_in[32]),
    .inData_33(stage_4_per_in[33]),
    .inData_34(stage_4_per_in[34]),
    .inData_35(stage_4_per_in[35]),
    .inData_36(stage_4_per_in[36]),
    .inData_37(stage_4_per_in[37]),
    .inData_38(stage_4_per_in[38]),
    .inData_39(stage_4_per_in[39]),
    .inData_40(stage_4_per_in[40]),
    .inData_41(stage_4_per_in[41]),
    .inData_42(stage_4_per_in[42]),
    .inData_43(stage_4_per_in[43]),
    .inData_44(stage_4_per_in[44]),
    .inData_45(stage_4_per_in[45]),
    .inData_46(stage_4_per_in[46]),
    .inData_47(stage_4_per_in[47]),
    .inData_48(stage_4_per_in[48]),
    .inData_49(stage_4_per_in[49]),
    .inData_50(stage_4_per_in[50]),
    .inData_51(stage_4_per_in[51]),
    .inData_52(stage_4_per_in[52]),
    .inData_53(stage_4_per_in[53]),
    .inData_54(stage_4_per_in[54]),
    .inData_55(stage_4_per_in[55]),
    .inData_56(stage_4_per_in[56]),
    .inData_57(stage_4_per_in[57]),
    .inData_58(stage_4_per_in[58]),
    .inData_59(stage_4_per_in[59]),
    .inData_60(stage_4_per_in[60]),
    .inData_61(stage_4_per_in[61]),
    .inData_62(stage_4_per_in[62]),
    .inData_63(stage_4_per_in[63]),
    .outData_0(stage_4_per_out[0]),
    .outData_1(stage_4_per_out[1]),
    .outData_2(stage_4_per_out[2]),
    .outData_3(stage_4_per_out[3]),
    .outData_4(stage_4_per_out[4]),
    .outData_5(stage_4_per_out[5]),
    .outData_6(stage_4_per_out[6]),
    .outData_7(stage_4_per_out[7]),
    .outData_8(stage_4_per_out[8]),
    .outData_9(stage_4_per_out[9]),
    .outData_10(stage_4_per_out[10]),
    .outData_11(stage_4_per_out[11]),
    .outData_12(stage_4_per_out[12]),
    .outData_13(stage_4_per_out[13]),
    .outData_14(stage_4_per_out[14]),
    .outData_15(stage_4_per_out[15]),
    .outData_16(stage_4_per_out[16]),
    .outData_17(stage_4_per_out[17]),
    .outData_18(stage_4_per_out[18]),
    .outData_19(stage_4_per_out[19]),
    .outData_20(stage_4_per_out[20]),
    .outData_21(stage_4_per_out[21]),
    .outData_22(stage_4_per_out[22]),
    .outData_23(stage_4_per_out[23]),
    .outData_24(stage_4_per_out[24]),
    .outData_25(stage_4_per_out[25]),
    .outData_26(stage_4_per_out[26]),
    .outData_27(stage_4_per_out[27]),
    .outData_28(stage_4_per_out[28]),
    .outData_29(stage_4_per_out[29]),
    .outData_30(stage_4_per_out[30]),
    .outData_31(stage_4_per_out[31]),
    .outData_32(stage_4_per_out[32]),
    .outData_33(stage_4_per_out[33]),
    .outData_34(stage_4_per_out[34]),
    .outData_35(stage_4_per_out[35]),
    .outData_36(stage_4_per_out[36]),
    .outData_37(stage_4_per_out[37]),
    .outData_38(stage_4_per_out[38]),
    .outData_39(stage_4_per_out[39]),
    .outData_40(stage_4_per_out[40]),
    .outData_41(stage_4_per_out[41]),
    .outData_42(stage_4_per_out[42]),
    .outData_43(stage_4_per_out[43]),
    .outData_44(stage_4_per_out[44]),
    .outData_45(stage_4_per_out[45]),
    .outData_46(stage_4_per_out[46]),
    .outData_47(stage_4_per_out[47]),
    .outData_48(stage_4_per_out[48]),
    .outData_49(stage_4_per_out[49]),
    .outData_50(stage_4_per_out[50]),
    .outData_51(stage_4_per_out[51]),
    .outData_52(stage_4_per_out[52]),
    .outData_53(stage_4_per_out[53]),
    .outData_54(stage_4_per_out[54]),
    .outData_55(stage_4_per_out[55]),
    .outData_56(stage_4_per_out[56]),
    .outData_57(stage_4_per_out[57]),
    .outData_58(stage_4_per_out[58]),
    .outData_59(stage_4_per_out[59]),
    .outData_60(stage_4_per_out[60]),
    .outData_61(stage_4_per_out[61]),
    .outData_62(stage_4_per_out[62]),
    .outData_63(stage_4_per_out[63]),
    .in_start(in_start[4]),
    .out_start(out_start[4]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 5 32 butterfly units
  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_0 (
    .x_in(stage_4_per_out[0]),
    .y_in(stage_4_per_out[1]),
    .x_out(stage_5_per_in[0]),
    .y_out(stage_5_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_1 (
    .x_in(stage_4_per_out[2]),
    .y_in(stage_4_per_out[3]),
    .x_out(stage_5_per_in[2]),
    .y_out(stage_5_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_2 (
    .x_in(stage_4_per_out[4]),
    .y_in(stage_4_per_out[5]),
    .x_out(stage_5_per_in[4]),
    .y_out(stage_5_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_3 (
    .x_in(stage_4_per_out[6]),
    .y_in(stage_4_per_out[7]),
    .x_out(stage_5_per_in[6]),
    .y_out(stage_5_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_4 (
    .x_in(stage_4_per_out[8]),
    .y_in(stage_4_per_out[9]),
    .x_out(stage_5_per_in[8]),
    .y_out(stage_5_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_5 (
    .x_in(stage_4_per_out[10]),
    .y_in(stage_4_per_out[11]),
    .x_out(stage_5_per_in[10]),
    .y_out(stage_5_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_6 (
    .x_in(stage_4_per_out[12]),
    .y_in(stage_4_per_out[13]),
    .x_out(stage_5_per_in[12]),
    .y_out(stage_5_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_7 (
    .x_in(stage_4_per_out[14]),
    .y_in(stage_4_per_out[15]),
    .x_out(stage_5_per_in[14]),
    .y_out(stage_5_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_8 (
    .x_in(stage_4_per_out[16]),
    .y_in(stage_4_per_out[17]),
    .x_out(stage_5_per_in[16]),
    .y_out(stage_5_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_9 (
    .x_in(stage_4_per_out[18]),
    .y_in(stage_4_per_out[19]),
    .x_out(stage_5_per_in[18]),
    .y_out(stage_5_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_10 (
    .x_in(stage_4_per_out[20]),
    .y_in(stage_4_per_out[21]),
    .x_out(stage_5_per_in[20]),
    .y_out(stage_5_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_11 (
    .x_in(stage_4_per_out[22]),
    .y_in(stage_4_per_out[23]),
    .x_out(stage_5_per_in[22]),
    .y_out(stage_5_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_12 (
    .x_in(stage_4_per_out[24]),
    .y_in(stage_4_per_out[25]),
    .x_out(stage_5_per_in[24]),
    .y_out(stage_5_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_13 (
    .x_in(stage_4_per_out[26]),
    .y_in(stage_4_per_out[27]),
    .x_out(stage_5_per_in[26]),
    .y_out(stage_5_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_14 (
    .x_in(stage_4_per_out[28]),
    .y_in(stage_4_per_out[29]),
    .x_out(stage_5_per_in[28]),
    .y_out(stage_5_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_15 (
    .x_in(stage_4_per_out[30]),
    .y_in(stage_4_per_out[31]),
    .x_out(stage_5_per_in[30]),
    .y_out(stage_5_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_16 (
    .x_in(stage_4_per_out[32]),
    .y_in(stage_4_per_out[33]),
    .x_out(stage_5_per_in[32]),
    .y_out(stage_5_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_17 (
    .x_in(stage_4_per_out[34]),
    .y_in(stage_4_per_out[35]),
    .x_out(stage_5_per_in[34]),
    .y_out(stage_5_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_18 (
    .x_in(stage_4_per_out[36]),
    .y_in(stage_4_per_out[37]),
    .x_out(stage_5_per_in[36]),
    .y_out(stage_5_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_19 (
    .x_in(stage_4_per_out[38]),
    .y_in(stage_4_per_out[39]),
    .x_out(stage_5_per_in[38]),
    .y_out(stage_5_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_20 (
    .x_in(stage_4_per_out[40]),
    .y_in(stage_4_per_out[41]),
    .x_out(stage_5_per_in[40]),
    .y_out(stage_5_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_21 (
    .x_in(stage_4_per_out[42]),
    .y_in(stage_4_per_out[43]),
    .x_out(stage_5_per_in[42]),
    .y_out(stage_5_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_22 (
    .x_in(stage_4_per_out[44]),
    .y_in(stage_4_per_out[45]),
    .x_out(stage_5_per_in[44]),
    .y_out(stage_5_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_23 (
    .x_in(stage_4_per_out[46]),
    .y_in(stage_4_per_out[47]),
    .x_out(stage_5_per_in[46]),
    .y_out(stage_5_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_24 (
    .x_in(stage_4_per_out[48]),
    .y_in(stage_4_per_out[49]),
    .x_out(stage_5_per_in[48]),
    .y_out(stage_5_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_25 (
    .x_in(stage_4_per_out[50]),
    .y_in(stage_4_per_out[51]),
    .x_out(stage_5_per_in[50]),
    .y_out(stage_5_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_26 (
    .x_in(stage_4_per_out[52]),
    .y_in(stage_4_per_out[53]),
    .x_out(stage_5_per_in[52]),
    .y_out(stage_5_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_27 (
    .x_in(stage_4_per_out[54]),
    .y_in(stage_4_per_out[55]),
    .x_out(stage_5_per_in[54]),
    .y_out(stage_5_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_28 (
    .x_in(stage_4_per_out[56]),
    .y_in(stage_4_per_out[57]),
    .x_out(stage_5_per_in[56]),
    .y_out(stage_5_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_29 (
    .x_in(stage_4_per_out[58]),
    .y_in(stage_4_per_out[59]),
    .x_out(stage_5_per_in[58]),
    .y_out(stage_5_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_30 (
    .x_in(stage_4_per_out[60]),
    .y_in(stage_4_per_out[61]),
    .x_out(stage_5_per_in[60]),
    .y_out(stage_5_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 185598009, 239095400, 39593842, 169276669, 141548072, 197386970, 119224607,
              159115155, 208403048, 102065274, 111284191, 157028693, 30748955, 210568560, 91114882,
              74680748, 162373432, 155896930, 145384235, 100099056, 71471012, 136571165, 33165861,
              149429971, 206324144, 175609590, 152865265, 201062854, 138074788, 191727270, 41084242,
              227611463, 196909902, 49823188, 78852289, 202366126, 146694818, 120670867, 86517113,
              256674305, 114407843, 233560477, 78462606, 92577793, 70582130, 172642311, 215696667,
              251290023, 193045667, 202257393, 242795574, 240684902, 47317233, 263678998, 152412548,
              200054106, 76707105, 140204941, 170752771, 109553202, 179817683, 262046585, 165226744}))
  stage_5_butterfly_31 (
    .x_in(stage_4_per_out[62]),
    .y_in(stage_4_per_out[63]),
    .x_out(stage_5_per_in[62]),
    .y_out(stage_5_per_in[63]),
    .clk(clk),
    .rst(rst)
  );



  // TODO(Yang): stage 5 -> stage 6 permutation
  // FIXME: ignore butterfly units for now.
  stage_5_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_5_6_per (
    .inData_0(stage_5_per_in[0]),
    .inData_1(stage_5_per_in[1]),
    .inData_2(stage_5_per_in[2]),
    .inData_3(stage_5_per_in[3]),
    .inData_4(stage_5_per_in[4]),
    .inData_5(stage_5_per_in[5]),
    .inData_6(stage_5_per_in[6]),
    .inData_7(stage_5_per_in[7]),
    .inData_8(stage_5_per_in[8]),
    .inData_9(stage_5_per_in[9]),
    .inData_10(stage_5_per_in[10]),
    .inData_11(stage_5_per_in[11]),
    .inData_12(stage_5_per_in[12]),
    .inData_13(stage_5_per_in[13]),
    .inData_14(stage_5_per_in[14]),
    .inData_15(stage_5_per_in[15]),
    .inData_16(stage_5_per_in[16]),
    .inData_17(stage_5_per_in[17]),
    .inData_18(stage_5_per_in[18]),
    .inData_19(stage_5_per_in[19]),
    .inData_20(stage_5_per_in[20]),
    .inData_21(stage_5_per_in[21]),
    .inData_22(stage_5_per_in[22]),
    .inData_23(stage_5_per_in[23]),
    .inData_24(stage_5_per_in[24]),
    .inData_25(stage_5_per_in[25]),
    .inData_26(stage_5_per_in[26]),
    .inData_27(stage_5_per_in[27]),
    .inData_28(stage_5_per_in[28]),
    .inData_29(stage_5_per_in[29]),
    .inData_30(stage_5_per_in[30]),
    .inData_31(stage_5_per_in[31]),
    .inData_32(stage_5_per_in[32]),
    .inData_33(stage_5_per_in[33]),
    .inData_34(stage_5_per_in[34]),
    .inData_35(stage_5_per_in[35]),
    .inData_36(stage_5_per_in[36]),
    .inData_37(stage_5_per_in[37]),
    .inData_38(stage_5_per_in[38]),
    .inData_39(stage_5_per_in[39]),
    .inData_40(stage_5_per_in[40]),
    .inData_41(stage_5_per_in[41]),
    .inData_42(stage_5_per_in[42]),
    .inData_43(stage_5_per_in[43]),
    .inData_44(stage_5_per_in[44]),
    .inData_45(stage_5_per_in[45]),
    .inData_46(stage_5_per_in[46]),
    .inData_47(stage_5_per_in[47]),
    .inData_48(stage_5_per_in[48]),
    .inData_49(stage_5_per_in[49]),
    .inData_50(stage_5_per_in[50]),
    .inData_51(stage_5_per_in[51]),
    .inData_52(stage_5_per_in[52]),
    .inData_53(stage_5_per_in[53]),
    .inData_54(stage_5_per_in[54]),
    .inData_55(stage_5_per_in[55]),
    .inData_56(stage_5_per_in[56]),
    .inData_57(stage_5_per_in[57]),
    .inData_58(stage_5_per_in[58]),
    .inData_59(stage_5_per_in[59]),
    .inData_60(stage_5_per_in[60]),
    .inData_61(stage_5_per_in[61]),
    .inData_62(stage_5_per_in[62]),
    .inData_63(stage_5_per_in[63]),
    .outData_0(stage_5_per_out[0]),
    .outData_1(stage_5_per_out[1]),
    .outData_2(stage_5_per_out[2]),
    .outData_3(stage_5_per_out[3]),
    .outData_4(stage_5_per_out[4]),
    .outData_5(stage_5_per_out[5]),
    .outData_6(stage_5_per_out[6]),
    .outData_7(stage_5_per_out[7]),
    .outData_8(stage_5_per_out[8]),
    .outData_9(stage_5_per_out[9]),
    .outData_10(stage_5_per_out[10]),
    .outData_11(stage_5_per_out[11]),
    .outData_12(stage_5_per_out[12]),
    .outData_13(stage_5_per_out[13]),
    .outData_14(stage_5_per_out[14]),
    .outData_15(stage_5_per_out[15]),
    .outData_16(stage_5_per_out[16]),
    .outData_17(stage_5_per_out[17]),
    .outData_18(stage_5_per_out[18]),
    .outData_19(stage_5_per_out[19]),
    .outData_20(stage_5_per_out[20]),
    .outData_21(stage_5_per_out[21]),
    .outData_22(stage_5_per_out[22]),
    .outData_23(stage_5_per_out[23]),
    .outData_24(stage_5_per_out[24]),
    .outData_25(stage_5_per_out[25]),
    .outData_26(stage_5_per_out[26]),
    .outData_27(stage_5_per_out[27]),
    .outData_28(stage_5_per_out[28]),
    .outData_29(stage_5_per_out[29]),
    .outData_30(stage_5_per_out[30]),
    .outData_31(stage_5_per_out[31]),
    .outData_32(stage_5_per_out[32]),
    .outData_33(stage_5_per_out[33]),
    .outData_34(stage_5_per_out[34]),
    .outData_35(stage_5_per_out[35]),
    .outData_36(stage_5_per_out[36]),
    .outData_37(stage_5_per_out[37]),
    .outData_38(stage_5_per_out[38]),
    .outData_39(stage_5_per_out[39]),
    .outData_40(stage_5_per_out[40]),
    .outData_41(stage_5_per_out[41]),
    .outData_42(stage_5_per_out[42]),
    .outData_43(stage_5_per_out[43]),
    .outData_44(stage_5_per_out[44]),
    .outData_45(stage_5_per_out[45]),
    .outData_46(stage_5_per_out[46]),
    .outData_47(stage_5_per_out[47]),
    .outData_48(stage_5_per_out[48]),
    .outData_49(stage_5_per_out[49]),
    .outData_50(stage_5_per_out[50]),
    .outData_51(stage_5_per_out[51]),
    .outData_52(stage_5_per_out[52]),
    .outData_53(stage_5_per_out[53]),
    .outData_54(stage_5_per_out[54]),
    .outData_55(stage_5_per_out[55]),
    .outData_56(stage_5_per_out[56]),
    .outData_57(stage_5_per_out[57]),
    .outData_58(stage_5_per_out[58]),
    .outData_59(stage_5_per_out[59]),
    .outData_60(stage_5_per_out[60]),
    .outData_61(stage_5_per_out[61]),
    .outData_62(stage_5_per_out[62]),
    .outData_63(stage_5_per_out[63]),
    .in_start(in_start[5]),
    .out_start(out_start[5]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 6 32 butterfly units
  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_0 (
    .x_in(stage_5_per_out[0]),
    .y_in(stage_5_per_out[1]),
    .x_out(stage_6_per_in[0]),
    .y_out(stage_6_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_1 (
    .x_in(stage_5_per_out[2]),
    .y_in(stage_5_per_out[3]),
    .x_out(stage_6_per_in[2]),
    .y_out(stage_6_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_2 (
    .x_in(stage_5_per_out[4]),
    .y_in(stage_5_per_out[5]),
    .x_out(stage_6_per_in[4]),
    .y_out(stage_6_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_3 (
    .x_in(stage_5_per_out[6]),
    .y_in(stage_5_per_out[7]),
    .x_out(stage_6_per_in[6]),
    .y_out(stage_6_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_4 (
    .x_in(stage_5_per_out[8]),
    .y_in(stage_5_per_out[9]),
    .x_out(stage_6_per_in[8]),
    .y_out(stage_6_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_5 (
    .x_in(stage_5_per_out[10]),
    .y_in(stage_5_per_out[11]),
    .x_out(stage_6_per_in[10]),
    .y_out(stage_6_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_6 (
    .x_in(stage_5_per_out[12]),
    .y_in(stage_5_per_out[13]),
    .x_out(stage_6_per_in[12]),
    .y_out(stage_6_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_7 (
    .x_in(stage_5_per_out[14]),
    .y_in(stage_5_per_out[15]),
    .x_out(stage_6_per_in[14]),
    .y_out(stage_6_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_8 (
    .x_in(stage_5_per_out[16]),
    .y_in(stage_5_per_out[17]),
    .x_out(stage_6_per_in[16]),
    .y_out(stage_6_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_9 (
    .x_in(stage_5_per_out[18]),
    .y_in(stage_5_per_out[19]),
    .x_out(stage_6_per_in[18]),
    .y_out(stage_6_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_10 (
    .x_in(stage_5_per_out[20]),
    .y_in(stage_5_per_out[21]),
    .x_out(stage_6_per_in[20]),
    .y_out(stage_6_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_11 (
    .x_in(stage_5_per_out[22]),
    .y_in(stage_5_per_out[23]),
    .x_out(stage_6_per_in[22]),
    .y_out(stage_6_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_12 (
    .x_in(stage_5_per_out[24]),
    .y_in(stage_5_per_out[25]),
    .x_out(stage_6_per_in[24]),
    .y_out(stage_6_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_13 (
    .x_in(stage_5_per_out[26]),
    .y_in(stage_5_per_out[27]),
    .x_out(stage_6_per_in[26]),
    .y_out(stage_6_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_14 (
    .x_in(stage_5_per_out[28]),
    .y_in(stage_5_per_out[29]),
    .x_out(stage_6_per_in[28]),
    .y_out(stage_6_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_15 (
    .x_in(stage_5_per_out[30]),
    .y_in(stage_5_per_out[31]),
    .x_out(stage_6_per_in[30]),
    .y_out(stage_6_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_16 (
    .x_in(stage_5_per_out[32]),
    .y_in(stage_5_per_out[33]),
    .x_out(stage_6_per_in[32]),
    .y_out(stage_6_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_17 (
    .x_in(stage_5_per_out[34]),
    .y_in(stage_5_per_out[35]),
    .x_out(stage_6_per_in[34]),
    .y_out(stage_6_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_18 (
    .x_in(stage_5_per_out[36]),
    .y_in(stage_5_per_out[37]),
    .x_out(stage_6_per_in[36]),
    .y_out(stage_6_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_19 (
    .x_in(stage_5_per_out[38]),
    .y_in(stage_5_per_out[39]),
    .x_out(stage_6_per_in[38]),
    .y_out(stage_6_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_20 (
    .x_in(stage_5_per_out[40]),
    .y_in(stage_5_per_out[41]),
    .x_out(stage_6_per_in[40]),
    .y_out(stage_6_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_21 (
    .x_in(stage_5_per_out[42]),
    .y_in(stage_5_per_out[43]),
    .x_out(stage_6_per_in[42]),
    .y_out(stage_6_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_22 (
    .x_in(stage_5_per_out[44]),
    .y_in(stage_5_per_out[45]),
    .x_out(stage_6_per_in[44]),
    .y_out(stage_6_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_23 (
    .x_in(stage_5_per_out[46]),
    .y_in(stage_5_per_out[47]),
    .x_out(stage_6_per_in[46]),
    .y_out(stage_6_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_24 (
    .x_in(stage_5_per_out[48]),
    .y_in(stage_5_per_out[49]),
    .x_out(stage_6_per_in[48]),
    .y_out(stage_6_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_25 (
    .x_in(stage_5_per_out[50]),
    .y_in(stage_5_per_out[51]),
    .x_out(stage_6_per_in[50]),
    .y_out(stage_6_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_26 (
    .x_in(stage_5_per_out[52]),
    .y_in(stage_5_per_out[53]),
    .x_out(stage_6_per_in[52]),
    .y_out(stage_6_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_27 (
    .x_in(stage_5_per_out[54]),
    .y_in(stage_5_per_out[55]),
    .x_out(stage_6_per_in[54]),
    .y_out(stage_6_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_28 (
    .x_in(stage_5_per_out[56]),
    .y_in(stage_5_per_out[57]),
    .x_out(stage_6_per_in[56]),
    .y_out(stage_6_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_29 (
    .x_in(stage_5_per_out[58]),
    .y_in(stage_5_per_out[59]),
    .x_out(stage_6_per_in[58]),
    .y_out(stage_6_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_30 (
    .x_in(stage_5_per_out[60]),
    .y_in(stage_5_per_out[61]),
    .x_out(stage_6_per_in[60]),
    .y_out(stage_6_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 102773617, 102773617, 210831626, 210831626, 84893967, 84893967,
              119480423, 119480423, 102579498, 102579498, 129001811, 129001811, 72061017, 72061017,
              72052889, 72052889, 73825164, 73825164, 18533839, 18533839, 168579404, 168579404,
              47877183, 47877183, 184798272, 184798272, 5258704, 5258704, 92744225, 92744225,
              221840088, 221840088, 216372172, 216372172, 231414272, 231414272, 94135184, 94135184,
              89995519, 89995519, 220656190, 220656190, 183300662, 183300662, 160020761, 160020761,
              249274747, 249274747, 62061822, 62061822, 76573097, 76573097, 35289455, 35289455,
              234642902, 234642902, 229105823, 229105823, 256670830, 256670830, 143639106, 143639106}))
  stage_6_butterfly_31 (
    .x_in(stage_5_per_out[62]),
    .y_in(stage_5_per_out[63]),
    .x_out(stage_6_per_in[62]),
    .y_out(stage_6_per_in[63]),
    .clk(clk),
    .rst(rst)
  );



  // TODO(Yang): stage 6 -> stage 7 permutation
  // FIXME: ignore butterfly units for now.
  stage_6_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_6_7_per (
    .inData_0(stage_6_per_in[0]),
    .inData_1(stage_6_per_in[1]),
    .inData_2(stage_6_per_in[2]),
    .inData_3(stage_6_per_in[3]),
    .inData_4(stage_6_per_in[4]),
    .inData_5(stage_6_per_in[5]),
    .inData_6(stage_6_per_in[6]),
    .inData_7(stage_6_per_in[7]),
    .inData_8(stage_6_per_in[8]),
    .inData_9(stage_6_per_in[9]),
    .inData_10(stage_6_per_in[10]),
    .inData_11(stage_6_per_in[11]),
    .inData_12(stage_6_per_in[12]),
    .inData_13(stage_6_per_in[13]),
    .inData_14(stage_6_per_in[14]),
    .inData_15(stage_6_per_in[15]),
    .inData_16(stage_6_per_in[16]),
    .inData_17(stage_6_per_in[17]),
    .inData_18(stage_6_per_in[18]),
    .inData_19(stage_6_per_in[19]),
    .inData_20(stage_6_per_in[20]),
    .inData_21(stage_6_per_in[21]),
    .inData_22(stage_6_per_in[22]),
    .inData_23(stage_6_per_in[23]),
    .inData_24(stage_6_per_in[24]),
    .inData_25(stage_6_per_in[25]),
    .inData_26(stage_6_per_in[26]),
    .inData_27(stage_6_per_in[27]),
    .inData_28(stage_6_per_in[28]),
    .inData_29(stage_6_per_in[29]),
    .inData_30(stage_6_per_in[30]),
    .inData_31(stage_6_per_in[31]),
    .inData_32(stage_6_per_in[32]),
    .inData_33(stage_6_per_in[33]),
    .inData_34(stage_6_per_in[34]),
    .inData_35(stage_6_per_in[35]),
    .inData_36(stage_6_per_in[36]),
    .inData_37(stage_6_per_in[37]),
    .inData_38(stage_6_per_in[38]),
    .inData_39(stage_6_per_in[39]),
    .inData_40(stage_6_per_in[40]),
    .inData_41(stage_6_per_in[41]),
    .inData_42(stage_6_per_in[42]),
    .inData_43(stage_6_per_in[43]),
    .inData_44(stage_6_per_in[44]),
    .inData_45(stage_6_per_in[45]),
    .inData_46(stage_6_per_in[46]),
    .inData_47(stage_6_per_in[47]),
    .inData_48(stage_6_per_in[48]),
    .inData_49(stage_6_per_in[49]),
    .inData_50(stage_6_per_in[50]),
    .inData_51(stage_6_per_in[51]),
    .inData_52(stage_6_per_in[52]),
    .inData_53(stage_6_per_in[53]),
    .inData_54(stage_6_per_in[54]),
    .inData_55(stage_6_per_in[55]),
    .inData_56(stage_6_per_in[56]),
    .inData_57(stage_6_per_in[57]),
    .inData_58(stage_6_per_in[58]),
    .inData_59(stage_6_per_in[59]),
    .inData_60(stage_6_per_in[60]),
    .inData_61(stage_6_per_in[61]),
    .inData_62(stage_6_per_in[62]),
    .inData_63(stage_6_per_in[63]),
    .outData_0(stage_6_per_out[0]),
    .outData_1(stage_6_per_out[1]),
    .outData_2(stage_6_per_out[2]),
    .outData_3(stage_6_per_out[3]),
    .outData_4(stage_6_per_out[4]),
    .outData_5(stage_6_per_out[5]),
    .outData_6(stage_6_per_out[6]),
    .outData_7(stage_6_per_out[7]),
    .outData_8(stage_6_per_out[8]),
    .outData_9(stage_6_per_out[9]),
    .outData_10(stage_6_per_out[10]),
    .outData_11(stage_6_per_out[11]),
    .outData_12(stage_6_per_out[12]),
    .outData_13(stage_6_per_out[13]),
    .outData_14(stage_6_per_out[14]),
    .outData_15(stage_6_per_out[15]),
    .outData_16(stage_6_per_out[16]),
    .outData_17(stage_6_per_out[17]),
    .outData_18(stage_6_per_out[18]),
    .outData_19(stage_6_per_out[19]),
    .outData_20(stage_6_per_out[20]),
    .outData_21(stage_6_per_out[21]),
    .outData_22(stage_6_per_out[22]),
    .outData_23(stage_6_per_out[23]),
    .outData_24(stage_6_per_out[24]),
    .outData_25(stage_6_per_out[25]),
    .outData_26(stage_6_per_out[26]),
    .outData_27(stage_6_per_out[27]),
    .outData_28(stage_6_per_out[28]),
    .outData_29(stage_6_per_out[29]),
    .outData_30(stage_6_per_out[30]),
    .outData_31(stage_6_per_out[31]),
    .outData_32(stage_6_per_out[32]),
    .outData_33(stage_6_per_out[33]),
    .outData_34(stage_6_per_out[34]),
    .outData_35(stage_6_per_out[35]),
    .outData_36(stage_6_per_out[36]),
    .outData_37(stage_6_per_out[37]),
    .outData_38(stage_6_per_out[38]),
    .outData_39(stage_6_per_out[39]),
    .outData_40(stage_6_per_out[40]),
    .outData_41(stage_6_per_out[41]),
    .outData_42(stage_6_per_out[42]),
    .outData_43(stage_6_per_out[43]),
    .outData_44(stage_6_per_out[44]),
    .outData_45(stage_6_per_out[45]),
    .outData_46(stage_6_per_out[46]),
    .outData_47(stage_6_per_out[47]),
    .outData_48(stage_6_per_out[48]),
    .outData_49(stage_6_per_out[49]),
    .outData_50(stage_6_per_out[50]),
    .outData_51(stage_6_per_out[51]),
    .outData_52(stage_6_per_out[52]),
    .outData_53(stage_6_per_out[53]),
    .outData_54(stage_6_per_out[54]),
    .outData_55(stage_6_per_out[55]),
    .outData_56(stage_6_per_out[56]),
    .outData_57(stage_6_per_out[57]),
    .outData_58(stage_6_per_out[58]),
    .outData_59(stage_6_per_out[59]),
    .outData_60(stage_6_per_out[60]),
    .outData_61(stage_6_per_out[61]),
    .outData_62(stage_6_per_out[62]),
    .outData_63(stage_6_per_out[63]),
    .in_start(in_start[6]),
    .out_start(out_start[6]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 7 32 butterfly units
  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_0 (
    .x_in(stage_6_per_out[0]),
    .y_in(stage_6_per_out[1]),
    .x_out(stage_7_per_in[0]),
    .y_out(stage_7_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_1 (
    .x_in(stage_6_per_out[2]),
    .y_in(stage_6_per_out[3]),
    .x_out(stage_7_per_in[2]),
    .y_out(stage_7_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_2 (
    .x_in(stage_6_per_out[4]),
    .y_in(stage_6_per_out[5]),
    .x_out(stage_7_per_in[4]),
    .y_out(stage_7_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_3 (
    .x_in(stage_6_per_out[6]),
    .y_in(stage_6_per_out[7]),
    .x_out(stage_7_per_in[6]),
    .y_out(stage_7_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_4 (
    .x_in(stage_6_per_out[8]),
    .y_in(stage_6_per_out[9]),
    .x_out(stage_7_per_in[8]),
    .y_out(stage_7_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_5 (
    .x_in(stage_6_per_out[10]),
    .y_in(stage_6_per_out[11]),
    .x_out(stage_7_per_in[10]),
    .y_out(stage_7_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_6 (
    .x_in(stage_6_per_out[12]),
    .y_in(stage_6_per_out[13]),
    .x_out(stage_7_per_in[12]),
    .y_out(stage_7_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_7 (
    .x_in(stage_6_per_out[14]),
    .y_in(stage_6_per_out[15]),
    .x_out(stage_7_per_in[14]),
    .y_out(stage_7_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_8 (
    .x_in(stage_6_per_out[16]),
    .y_in(stage_6_per_out[17]),
    .x_out(stage_7_per_in[16]),
    .y_out(stage_7_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_9 (
    .x_in(stage_6_per_out[18]),
    .y_in(stage_6_per_out[19]),
    .x_out(stage_7_per_in[18]),
    .y_out(stage_7_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_10 (
    .x_in(stage_6_per_out[20]),
    .y_in(stage_6_per_out[21]),
    .x_out(stage_7_per_in[20]),
    .y_out(stage_7_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_11 (
    .x_in(stage_6_per_out[22]),
    .y_in(stage_6_per_out[23]),
    .x_out(stage_7_per_in[22]),
    .y_out(stage_7_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_12 (
    .x_in(stage_6_per_out[24]),
    .y_in(stage_6_per_out[25]),
    .x_out(stage_7_per_in[24]),
    .y_out(stage_7_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_13 (
    .x_in(stage_6_per_out[26]),
    .y_in(stage_6_per_out[27]),
    .x_out(stage_7_per_in[26]),
    .y_out(stage_7_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_14 (
    .x_in(stage_6_per_out[28]),
    .y_in(stage_6_per_out[29]),
    .x_out(stage_7_per_in[28]),
    .y_out(stage_7_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_15 (
    .x_in(stage_6_per_out[30]),
    .y_in(stage_6_per_out[31]),
    .x_out(stage_7_per_in[30]),
    .y_out(stage_7_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_16 (
    .x_in(stage_6_per_out[32]),
    .y_in(stage_6_per_out[33]),
    .x_out(stage_7_per_in[32]),
    .y_out(stage_7_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_17 (
    .x_in(stage_6_per_out[34]),
    .y_in(stage_6_per_out[35]),
    .x_out(stage_7_per_in[34]),
    .y_out(stage_7_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_18 (
    .x_in(stage_6_per_out[36]),
    .y_in(stage_6_per_out[37]),
    .x_out(stage_7_per_in[36]),
    .y_out(stage_7_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_19 (
    .x_in(stage_6_per_out[38]),
    .y_in(stage_6_per_out[39]),
    .x_out(stage_7_per_in[38]),
    .y_out(stage_7_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_20 (
    .x_in(stage_6_per_out[40]),
    .y_in(stage_6_per_out[41]),
    .x_out(stage_7_per_in[40]),
    .y_out(stage_7_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_21 (
    .x_in(stage_6_per_out[42]),
    .y_in(stage_6_per_out[43]),
    .x_out(stage_7_per_in[42]),
    .y_out(stage_7_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_22 (
    .x_in(stage_6_per_out[44]),
    .y_in(stage_6_per_out[45]),
    .x_out(stage_7_per_in[44]),
    .y_out(stage_7_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_23 (
    .x_in(stage_6_per_out[46]),
    .y_in(stage_6_per_out[47]),
    .x_out(stage_7_per_in[46]),
    .y_out(stage_7_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_24 (
    .x_in(stage_6_per_out[48]),
    .y_in(stage_6_per_out[49]),
    .x_out(stage_7_per_in[48]),
    .y_out(stage_7_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_25 (
    .x_in(stage_6_per_out[50]),
    .y_in(stage_6_per_out[51]),
    .x_out(stage_7_per_in[50]),
    .y_out(stage_7_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_26 (
    .x_in(stage_6_per_out[52]),
    .y_in(stage_6_per_out[53]),
    .x_out(stage_7_per_in[52]),
    .y_out(stage_7_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_27 (
    .x_in(stage_6_per_out[54]),
    .y_in(stage_6_per_out[55]),
    .x_out(stage_7_per_in[54]),
    .y_out(stage_7_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_28 (
    .x_in(stage_6_per_out[56]),
    .y_in(stage_6_per_out[57]),
    .x_out(stage_7_per_in[56]),
    .y_out(stage_7_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_29 (
    .x_in(stage_6_per_out[58]),
    .y_in(stage_6_per_out[59]),
    .x_out(stage_7_per_in[58]),
    .y_out(stage_7_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_30 (
    .x_in(stage_6_per_out[60]),
    .y_in(stage_6_per_out[61]),
    .x_out(stage_7_per_in[60]),
    .y_out(stage_7_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_31 (
    .x_in(stage_6_per_out[62]),
    .y_in(stage_6_per_out[63]),
    .x_out(stage_7_per_in[62]),
    .y_out(stage_7_per_in[63]),
    .clk(clk),
    .rst(rst)
  );




  // TODO(Yang): stage 7 -> stage 8 permutation
  // FIXME: ignore butterfly units for now.
  stage_7_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_7_8_per (
    .inData_0(stage_7_per_in[0]),
    .inData_1(stage_7_per_in[1]),
    .inData_2(stage_7_per_in[2]),
    .inData_3(stage_7_per_in[3]),
    .inData_4(stage_7_per_in[4]),
    .inData_5(stage_7_per_in[5]),
    .inData_6(stage_7_per_in[6]),
    .inData_7(stage_7_per_in[7]),
    .inData_8(stage_7_per_in[8]),
    .inData_9(stage_7_per_in[9]),
    .inData_10(stage_7_per_in[10]),
    .inData_11(stage_7_per_in[11]),
    .inData_12(stage_7_per_in[12]),
    .inData_13(stage_7_per_in[13]),
    .inData_14(stage_7_per_in[14]),
    .inData_15(stage_7_per_in[15]),
    .inData_16(stage_7_per_in[16]),
    .inData_17(stage_7_per_in[17]),
    .inData_18(stage_7_per_in[18]),
    .inData_19(stage_7_per_in[19]),
    .inData_20(stage_7_per_in[20]),
    .inData_21(stage_7_per_in[21]),
    .inData_22(stage_7_per_in[22]),
    .inData_23(stage_7_per_in[23]),
    .inData_24(stage_7_per_in[24]),
    .inData_25(stage_7_per_in[25]),
    .inData_26(stage_7_per_in[26]),
    .inData_27(stage_7_per_in[27]),
    .inData_28(stage_7_per_in[28]),
    .inData_29(stage_7_per_in[29]),
    .inData_30(stage_7_per_in[30]),
    .inData_31(stage_7_per_in[31]),
    .inData_32(stage_7_per_in[32]),
    .inData_33(stage_7_per_in[33]),
    .inData_34(stage_7_per_in[34]),
    .inData_35(stage_7_per_in[35]),
    .inData_36(stage_7_per_in[36]),
    .inData_37(stage_7_per_in[37]),
    .inData_38(stage_7_per_in[38]),
    .inData_39(stage_7_per_in[39]),
    .inData_40(stage_7_per_in[40]),
    .inData_41(stage_7_per_in[41]),
    .inData_42(stage_7_per_in[42]),
    .inData_43(stage_7_per_in[43]),
    .inData_44(stage_7_per_in[44]),
    .inData_45(stage_7_per_in[45]),
    .inData_46(stage_7_per_in[46]),
    .inData_47(stage_7_per_in[47]),
    .inData_48(stage_7_per_in[48]),
    .inData_49(stage_7_per_in[49]),
    .inData_50(stage_7_per_in[50]),
    .inData_51(stage_7_per_in[51]),
    .inData_52(stage_7_per_in[52]),
    .inData_53(stage_7_per_in[53]),
    .inData_54(stage_7_per_in[54]),
    .inData_55(stage_7_per_in[55]),
    .inData_56(stage_7_per_in[56]),
    .inData_57(stage_7_per_in[57]),
    .inData_58(stage_7_per_in[58]),
    .inData_59(stage_7_per_in[59]),
    .inData_60(stage_7_per_in[60]),
    .inData_61(stage_7_per_in[61]),
    .inData_62(stage_7_per_in[62]),
    .inData_63(stage_7_per_in[63]),
    .outData_0(stage_7_per_out[0]),
    .outData_1(stage_7_per_out[1]),
    .outData_2(stage_7_per_out[2]),
    .outData_3(stage_7_per_out[3]),
    .outData_4(stage_7_per_out[4]),
    .outData_5(stage_7_per_out[5]),
    .outData_6(stage_7_per_out[6]),
    .outData_7(stage_7_per_out[7]),
    .outData_8(stage_7_per_out[8]),
    .outData_9(stage_7_per_out[9]),
    .outData_10(stage_7_per_out[10]),
    .outData_11(stage_7_per_out[11]),
    .outData_12(stage_7_per_out[12]),
    .outData_13(stage_7_per_out[13]),
    .outData_14(stage_7_per_out[14]),
    .outData_15(stage_7_per_out[15]),
    .outData_16(stage_7_per_out[16]),
    .outData_17(stage_7_per_out[17]),
    .outData_18(stage_7_per_out[18]),
    .outData_19(stage_7_per_out[19]),
    .outData_20(stage_7_per_out[20]),
    .outData_21(stage_7_per_out[21]),
    .outData_22(stage_7_per_out[22]),
    .outData_23(stage_7_per_out[23]),
    .outData_24(stage_7_per_out[24]),
    .outData_25(stage_7_per_out[25]),
    .outData_26(stage_7_per_out[26]),
    .outData_27(stage_7_per_out[27]),
    .outData_28(stage_7_per_out[28]),
    .outData_29(stage_7_per_out[29]),
    .outData_30(stage_7_per_out[30]),
    .outData_31(stage_7_per_out[31]),
    .outData_32(stage_7_per_out[32]),
    .outData_33(stage_7_per_out[33]),
    .outData_34(stage_7_per_out[34]),
    .outData_35(stage_7_per_out[35]),
    .outData_36(stage_7_per_out[36]),
    .outData_37(stage_7_per_out[37]),
    .outData_38(stage_7_per_out[38]),
    .outData_39(stage_7_per_out[39]),
    .outData_40(stage_7_per_out[40]),
    .outData_41(stage_7_per_out[41]),
    .outData_42(stage_7_per_out[42]),
    .outData_43(stage_7_per_out[43]),
    .outData_44(stage_7_per_out[44]),
    .outData_45(stage_7_per_out[45]),
    .outData_46(stage_7_per_out[46]),
    .outData_47(stage_7_per_out[47]),
    .outData_48(stage_7_per_out[48]),
    .outData_49(stage_7_per_out[49]),
    .outData_50(stage_7_per_out[50]),
    .outData_51(stage_7_per_out[51]),
    .outData_52(stage_7_per_out[52]),
    .outData_53(stage_7_per_out[53]),
    .outData_54(stage_7_per_out[54]),
    .outData_55(stage_7_per_out[55]),
    .outData_56(stage_7_per_out[56]),
    .outData_57(stage_7_per_out[57]),
    .outData_58(stage_7_per_out[58]),
    .outData_59(stage_7_per_out[59]),
    .outData_60(stage_7_per_out[60]),
    .outData_61(stage_7_per_out[61]),
    .outData_62(stage_7_per_out[62]),
    .outData_63(stage_7_per_out[63]),
    .in_start(in_start[7]),
    .out_start(out_start[7]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 8 32 butterfly units
  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_0 (
    .x_in(stage_7_per_out[0]),
    .y_in(stage_7_per_out[1]),
    .x_out(stage_8_per_in[0]),
    .y_out(stage_8_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_1 (
    .x_in(stage_7_per_out[2]),
    .y_in(stage_7_per_out[3]),
    .x_out(stage_8_per_in[2]),
    .y_out(stage_8_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_2 (
    .x_in(stage_7_per_out[4]),
    .y_in(stage_7_per_out[5]),
    .x_out(stage_8_per_in[4]),
    .y_out(stage_8_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_3 (
    .x_in(stage_7_per_out[6]),
    .y_in(stage_7_per_out[7]),
    .x_out(stage_8_per_in[6]),
    .y_out(stage_8_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_4 (
    .x_in(stage_7_per_out[8]),
    .y_in(stage_7_per_out[9]),
    .x_out(stage_8_per_in[8]),
    .y_out(stage_8_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_5 (
    .x_in(stage_7_per_out[10]),
    .y_in(stage_7_per_out[11]),
    .x_out(stage_8_per_in[10]),
    .y_out(stage_8_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_6 (
    .x_in(stage_7_per_out[12]),
    .y_in(stage_7_per_out[13]),
    .x_out(stage_8_per_in[12]),
    .y_out(stage_8_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_7 (
    .x_in(stage_7_per_out[14]),
    .y_in(stage_7_per_out[15]),
    .x_out(stage_8_per_in[14]),
    .y_out(stage_8_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_8 (
    .x_in(stage_7_per_out[16]),
    .y_in(stage_7_per_out[17]),
    .x_out(stage_8_per_in[16]),
    .y_out(stage_8_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_9 (
    .x_in(stage_7_per_out[18]),
    .y_in(stage_7_per_out[19]),
    .x_out(stage_8_per_in[18]),
    .y_out(stage_8_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_10 (
    .x_in(stage_7_per_out[20]),
    .y_in(stage_7_per_out[21]),
    .x_out(stage_8_per_in[20]),
    .y_out(stage_8_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_11 (
    .x_in(stage_7_per_out[22]),
    .y_in(stage_7_per_out[23]),
    .x_out(stage_8_per_in[22]),
    .y_out(stage_8_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_12 (
    .x_in(stage_7_per_out[24]),
    .y_in(stage_7_per_out[25]),
    .x_out(stage_8_per_in[24]),
    .y_out(stage_8_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_13 (
    .x_in(stage_7_per_out[26]),
    .y_in(stage_7_per_out[27]),
    .x_out(stage_8_per_in[26]),
    .y_out(stage_8_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_14 (
    .x_in(stage_7_per_out[28]),
    .y_in(stage_7_per_out[29]),
    .x_out(stage_8_per_in[28]),
    .y_out(stage_8_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_15 (
    .x_in(stage_7_per_out[30]),
    .y_in(stage_7_per_out[31]),
    .x_out(stage_8_per_in[30]),
    .y_out(stage_8_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_16 (
    .x_in(stage_7_per_out[32]),
    .y_in(stage_7_per_out[33]),
    .x_out(stage_8_per_in[32]),
    .y_out(stage_8_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_17 (
    .x_in(stage_7_per_out[34]),
    .y_in(stage_7_per_out[35]),
    .x_out(stage_8_per_in[34]),
    .y_out(stage_8_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_18 (
    .x_in(stage_7_per_out[36]),
    .y_in(stage_7_per_out[37]),
    .x_out(stage_8_per_in[36]),
    .y_out(stage_8_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_19 (
    .x_in(stage_7_per_out[38]),
    .y_in(stage_7_per_out[39]),
    .x_out(stage_8_per_in[38]),
    .y_out(stage_8_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_20 (
    .x_in(stage_7_per_out[40]),
    .y_in(stage_7_per_out[41]),
    .x_out(stage_8_per_in[40]),
    .y_out(stage_8_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_21 (
    .x_in(stage_7_per_out[42]),
    .y_in(stage_7_per_out[43]),
    .x_out(stage_8_per_in[42]),
    .y_out(stage_8_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_22 (
    .x_in(stage_7_per_out[44]),
    .y_in(stage_7_per_out[45]),
    .x_out(stage_8_per_in[44]),
    .y_out(stage_8_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_23 (
    .x_in(stage_7_per_out[46]),
    .y_in(stage_7_per_out[47]),
    .x_out(stage_8_per_in[46]),
    .y_out(stage_8_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_24 (
    .x_in(stage_7_per_out[48]),
    .y_in(stage_7_per_out[49]),
    .x_out(stage_8_per_in[48]),
    .y_out(stage_8_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_25 (
    .x_in(stage_7_per_out[50]),
    .y_in(stage_7_per_out[51]),
    .x_out(stage_8_per_in[50]),
    .y_out(stage_8_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_26 (
    .x_in(stage_7_per_out[52]),
    .y_in(stage_7_per_out[53]),
    .x_out(stage_8_per_in[52]),
    .y_out(stage_8_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_27 (
    .x_in(stage_7_per_out[54]),
    .y_in(stage_7_per_out[55]),
    .x_out(stage_8_per_in[54]),
    .y_out(stage_8_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_28 (
    .x_in(stage_7_per_out[56]),
    .y_in(stage_7_per_out[57]),
    .x_out(stage_8_per_in[56]),
    .y_out(stage_8_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_29 (
    .x_in(stage_7_per_out[58]),
    .y_in(stage_7_per_out[59]),
    .x_out(stage_8_per_in[58]),
    .y_out(stage_8_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_30 (
    .x_in(stage_7_per_out[60]),
    .y_in(stage_7_per_out[61]),
    .x_out(stage_8_per_in[60]),
    .y_out(stage_8_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_31 (
    .x_in(stage_7_per_out[62]),
    .y_in(stage_7_per_out[63]),
    .x_out(stage_8_per_in[62]),
    .y_out(stage_8_per_in[63]),
    .clk(clk),
    .rst(rst)
  );




  // TODO(Yang): stage 8 -> stage 9 permutation
  // FIXME: ignore butterfly units for now.
  stage_8_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_8_9_per (
    .inData_0(stage_8_per_in[0]),
    .inData_1(stage_8_per_in[1]),
    .inData_2(stage_8_per_in[2]),
    .inData_3(stage_8_per_in[3]),
    .inData_4(stage_8_per_in[4]),
    .inData_5(stage_8_per_in[5]),
    .inData_6(stage_8_per_in[6]),
    .inData_7(stage_8_per_in[7]),
    .inData_8(stage_8_per_in[8]),
    .inData_9(stage_8_per_in[9]),
    .inData_10(stage_8_per_in[10]),
    .inData_11(stage_8_per_in[11]),
    .inData_12(stage_8_per_in[12]),
    .inData_13(stage_8_per_in[13]),
    .inData_14(stage_8_per_in[14]),
    .inData_15(stage_8_per_in[15]),
    .inData_16(stage_8_per_in[16]),
    .inData_17(stage_8_per_in[17]),
    .inData_18(stage_8_per_in[18]),
    .inData_19(stage_8_per_in[19]),
    .inData_20(stage_8_per_in[20]),
    .inData_21(stage_8_per_in[21]),
    .inData_22(stage_8_per_in[22]),
    .inData_23(stage_8_per_in[23]),
    .inData_24(stage_8_per_in[24]),
    .inData_25(stage_8_per_in[25]),
    .inData_26(stage_8_per_in[26]),
    .inData_27(stage_8_per_in[27]),
    .inData_28(stage_8_per_in[28]),
    .inData_29(stage_8_per_in[29]),
    .inData_30(stage_8_per_in[30]),
    .inData_31(stage_8_per_in[31]),
    .inData_32(stage_8_per_in[32]),
    .inData_33(stage_8_per_in[33]),
    .inData_34(stage_8_per_in[34]),
    .inData_35(stage_8_per_in[35]),
    .inData_36(stage_8_per_in[36]),
    .inData_37(stage_8_per_in[37]),
    .inData_38(stage_8_per_in[38]),
    .inData_39(stage_8_per_in[39]),
    .inData_40(stage_8_per_in[40]),
    .inData_41(stage_8_per_in[41]),
    .inData_42(stage_8_per_in[42]),
    .inData_43(stage_8_per_in[43]),
    .inData_44(stage_8_per_in[44]),
    .inData_45(stage_8_per_in[45]),
    .inData_46(stage_8_per_in[46]),
    .inData_47(stage_8_per_in[47]),
    .inData_48(stage_8_per_in[48]),
    .inData_49(stage_8_per_in[49]),
    .inData_50(stage_8_per_in[50]),
    .inData_51(stage_8_per_in[51]),
    .inData_52(stage_8_per_in[52]),
    .inData_53(stage_8_per_in[53]),
    .inData_54(stage_8_per_in[54]),
    .inData_55(stage_8_per_in[55]),
    .inData_56(stage_8_per_in[56]),
    .inData_57(stage_8_per_in[57]),
    .inData_58(stage_8_per_in[58]),
    .inData_59(stage_8_per_in[59]),
    .inData_60(stage_8_per_in[60]),
    .inData_61(stage_8_per_in[61]),
    .inData_62(stage_8_per_in[62]),
    .inData_63(stage_8_per_in[63]),
    .outData_0(stage_8_per_out[0]),
    .outData_1(stage_8_per_out[1]),
    .outData_2(stage_8_per_out[2]),
    .outData_3(stage_8_per_out[3]),
    .outData_4(stage_8_per_out[4]),
    .outData_5(stage_8_per_out[5]),
    .outData_6(stage_8_per_out[6]),
    .outData_7(stage_8_per_out[7]),
    .outData_8(stage_8_per_out[8]),
    .outData_9(stage_8_per_out[9]),
    .outData_10(stage_8_per_out[10]),
    .outData_11(stage_8_per_out[11]),
    .outData_12(stage_8_per_out[12]),
    .outData_13(stage_8_per_out[13]),
    .outData_14(stage_8_per_out[14]),
    .outData_15(stage_8_per_out[15]),
    .outData_16(stage_8_per_out[16]),
    .outData_17(stage_8_per_out[17]),
    .outData_18(stage_8_per_out[18]),
    .outData_19(stage_8_per_out[19]),
    .outData_20(stage_8_per_out[20]),
    .outData_21(stage_8_per_out[21]),
    .outData_22(stage_8_per_out[22]),
    .outData_23(stage_8_per_out[23]),
    .outData_24(stage_8_per_out[24]),
    .outData_25(stage_8_per_out[25]),
    .outData_26(stage_8_per_out[26]),
    .outData_27(stage_8_per_out[27]),
    .outData_28(stage_8_per_out[28]),
    .outData_29(stage_8_per_out[29]),
    .outData_30(stage_8_per_out[30]),
    .outData_31(stage_8_per_out[31]),
    .outData_32(stage_8_per_out[32]),
    .outData_33(stage_8_per_out[33]),
    .outData_34(stage_8_per_out[34]),
    .outData_35(stage_8_per_out[35]),
    .outData_36(stage_8_per_out[36]),
    .outData_37(stage_8_per_out[37]),
    .outData_38(stage_8_per_out[38]),
    .outData_39(stage_8_per_out[39]),
    .outData_40(stage_8_per_out[40]),
    .outData_41(stage_8_per_out[41]),
    .outData_42(stage_8_per_out[42]),
    .outData_43(stage_8_per_out[43]),
    .outData_44(stage_8_per_out[44]),
    .outData_45(stage_8_per_out[45]),
    .outData_46(stage_8_per_out[46]),
    .outData_47(stage_8_per_out[47]),
    .outData_48(stage_8_per_out[48]),
    .outData_49(stage_8_per_out[49]),
    .outData_50(stage_8_per_out[50]),
    .outData_51(stage_8_per_out[51]),
    .outData_52(stage_8_per_out[52]),
    .outData_53(stage_8_per_out[53]),
    .outData_54(stage_8_per_out[54]),
    .outData_55(stage_8_per_out[55]),
    .outData_56(stage_8_per_out[56]),
    .outData_57(stage_8_per_out[57]),
    .outData_58(stage_8_per_out[58]),
    .outData_59(stage_8_per_out[59]),
    .outData_60(stage_8_per_out[60]),
    .outData_61(stage_8_per_out[61]),
    .outData_62(stage_8_per_out[62]),
    .outData_63(stage_8_per_out[63]),
    .in_start(in_start[8]),
    .out_start(out_start[8]),
    .clk(clk),
    .rst(rst)
  );

  // TODO(Tian): stage 9 32 butterfly units
  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_0 (
    .x_in(stage_8_per_out[0]),
    .y_in(stage_8_per_out[1]),
    .x_out(stage_9_per_in[0]),
    .y_out(stage_9_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_1 (
    .x_in(stage_8_per_out[2]),
    .y_in(stage_8_per_out[3]),
    .x_out(stage_9_per_in[2]),
    .y_out(stage_9_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_2 (
    .x_in(stage_8_per_out[4]),
    .y_in(stage_8_per_out[5]),
    .x_out(stage_9_per_in[4]),
    .y_out(stage_9_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_3 (
    .x_in(stage_8_per_out[6]),
    .y_in(stage_8_per_out[7]),
    .x_out(stage_9_per_in[6]),
    .y_out(stage_9_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_4 (
    .x_in(stage_8_per_out[8]),
    .y_in(stage_8_per_out[9]),
    .x_out(stage_9_per_in[8]),
    .y_out(stage_9_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_5 (
    .x_in(stage_8_per_out[10]),
    .y_in(stage_8_per_out[11]),
    .x_out(stage_9_per_in[10]),
    .y_out(stage_9_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_6 (
    .x_in(stage_8_per_out[12]),
    .y_in(stage_8_per_out[13]),
    .x_out(stage_9_per_in[12]),
    .y_out(stage_9_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_7 (
    .x_in(stage_8_per_out[14]),
    .y_in(stage_8_per_out[15]),
    .x_out(stage_9_per_in[14]),
    .y_out(stage_9_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_8 (
    .x_in(stage_8_per_out[16]),
    .y_in(stage_8_per_out[17]),
    .x_out(stage_9_per_in[16]),
    .y_out(stage_9_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_9 (
    .x_in(stage_8_per_out[18]),
    .y_in(stage_8_per_out[19]),
    .x_out(stage_9_per_in[18]),
    .y_out(stage_9_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_10 (
    .x_in(stage_8_per_out[20]),
    .y_in(stage_8_per_out[21]),
    .x_out(stage_9_per_in[20]),
    .y_out(stage_9_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_11 (
    .x_in(stage_8_per_out[22]),
    .y_in(stage_8_per_out[23]),
    .x_out(stage_9_per_in[22]),
    .y_out(stage_9_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_12 (
    .x_in(stage_8_per_out[24]),
    .y_in(stage_8_per_out[25]),
    .x_out(stage_9_per_in[24]),
    .y_out(stage_9_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_13 (
    .x_in(stage_8_per_out[26]),
    .y_in(stage_8_per_out[27]),
    .x_out(stage_9_per_in[26]),
    .y_out(stage_9_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_14 (
    .x_in(stage_8_per_out[28]),
    .y_in(stage_8_per_out[29]),
    .x_out(stage_9_per_in[28]),
    .y_out(stage_9_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_15 (
    .x_in(stage_8_per_out[30]),
    .y_in(stage_8_per_out[31]),
    .x_out(stage_9_per_in[30]),
    .y_out(stage_9_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_16 (
    .x_in(stage_8_per_out[32]),
    .y_in(stage_8_per_out[33]),
    .x_out(stage_9_per_in[32]),
    .y_out(stage_9_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_17 (
    .x_in(stage_8_per_out[34]),
    .y_in(stage_8_per_out[35]),
    .x_out(stage_9_per_in[34]),
    .y_out(stage_9_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_18 (
    .x_in(stage_8_per_out[36]),
    .y_in(stage_8_per_out[37]),
    .x_out(stage_9_per_in[36]),
    .y_out(stage_9_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_19 (
    .x_in(stage_8_per_out[38]),
    .y_in(stage_8_per_out[39]),
    .x_out(stage_9_per_in[38]),
    .y_out(stage_9_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_20 (
    .x_in(stage_8_per_out[40]),
    .y_in(stage_8_per_out[41]),
    .x_out(stage_9_per_in[40]),
    .y_out(stage_9_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_21 (
    .x_in(stage_8_per_out[42]),
    .y_in(stage_8_per_out[43]),
    .x_out(stage_9_per_in[42]),
    .y_out(stage_9_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_22 (
    .x_in(stage_8_per_out[44]),
    .y_in(stage_8_per_out[45]),
    .x_out(stage_9_per_in[44]),
    .y_out(stage_9_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_23 (
    .x_in(stage_8_per_out[46]),
    .y_in(stage_8_per_out[47]),
    .x_out(stage_9_per_in[46]),
    .y_out(stage_9_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_24 (
    .x_in(stage_8_per_out[48]),
    .y_in(stage_8_per_out[49]),
    .x_out(stage_9_per_in[48]),
    .y_out(stage_9_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_25 (
    .x_in(stage_8_per_out[50]),
    .y_in(stage_8_per_out[51]),
    .x_out(stage_9_per_in[50]),
    .y_out(stage_9_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_26 (
    .x_in(stage_8_per_out[52]),
    .y_in(stage_8_per_out[53]),
    .x_out(stage_9_per_in[52]),
    .y_out(stage_9_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_27 (
    .x_in(stage_8_per_out[54]),
    .y_in(stage_8_per_out[55]),
    .x_out(stage_9_per_in[54]),
    .y_out(stage_9_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_28 (
    .x_in(stage_8_per_out[56]),
    .y_in(stage_8_per_out[57]),
    .x_out(stage_9_per_in[56]),
    .y_out(stage_9_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_29 (
    .x_in(stage_8_per_out[58]),
    .y_in(stage_8_per_out[59]),
    .x_out(stage_9_per_in[58]),
    .y_out(stage_9_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_30 (
    .x_in(stage_8_per_out[60]),
    .y_in(stage_8_per_out[61]),
    .x_out(stage_9_per_in[60]),
    .y_out(stage_9_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_31 (
    .x_in(stage_8_per_out[62]),
    .y_in(stage_8_per_out[63]),
    .x_out(stage_9_per_in[62]),
    .y_out(stage_9_per_in[63]),
    .clk(clk),
    .rst(rst)
  );



  // TODO(Yang): stage 8 -> stage 9 permutation
  // FIXME: ignore butterfly units for now.
  stage_9_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_9_10_per (
    .inData_0(stage_9_per_in[0]),
    .inData_1(stage_9_per_in[1]),
    .inData_2(stage_9_per_in[2]),
    .inData_3(stage_9_per_in[3]),
    .inData_4(stage_9_per_in[4]),
    .inData_5(stage_9_per_in[5]),
    .inData_6(stage_9_per_in[6]),
    .inData_7(stage_9_per_in[7]),
    .inData_8(stage_9_per_in[8]),
    .inData_9(stage_9_per_in[9]),
    .inData_10(stage_9_per_in[10]),
    .inData_11(stage_9_per_in[11]),
    .inData_12(stage_9_per_in[12]),
    .inData_13(stage_9_per_in[13]),
    .inData_14(stage_9_per_in[14]),
    .inData_15(stage_9_per_in[15]),
    .inData_16(stage_9_per_in[16]),
    .inData_17(stage_9_per_in[17]),
    .inData_18(stage_9_per_in[18]),
    .inData_19(stage_9_per_in[19]),
    .inData_20(stage_9_per_in[20]),
    .inData_21(stage_9_per_in[21]),
    .inData_22(stage_9_per_in[22]),
    .inData_23(stage_9_per_in[23]),
    .inData_24(stage_9_per_in[24]),
    .inData_25(stage_9_per_in[25]),
    .inData_26(stage_9_per_in[26]),
    .inData_27(stage_9_per_in[27]),
    .inData_28(stage_9_per_in[28]),
    .inData_29(stage_9_per_in[29]),
    .inData_30(stage_9_per_in[30]),
    .inData_31(stage_9_per_in[31]),
    .inData_32(stage_9_per_in[32]),
    .inData_33(stage_9_per_in[33]),
    .inData_34(stage_9_per_in[34]),
    .inData_35(stage_9_per_in[35]),
    .inData_36(stage_9_per_in[36]),
    .inData_37(stage_9_per_in[37]),
    .inData_38(stage_9_per_in[38]),
    .inData_39(stage_9_per_in[39]),
    .inData_40(stage_9_per_in[40]),
    .inData_41(stage_9_per_in[41]),
    .inData_42(stage_9_per_in[42]),
    .inData_43(stage_9_per_in[43]),
    .inData_44(stage_9_per_in[44]),
    .inData_45(stage_9_per_in[45]),
    .inData_46(stage_9_per_in[46]),
    .inData_47(stage_9_per_in[47]),
    .inData_48(stage_9_per_in[48]),
    .inData_49(stage_9_per_in[49]),
    .inData_50(stage_9_per_in[50]),
    .inData_51(stage_9_per_in[51]),
    .inData_52(stage_9_per_in[52]),
    .inData_53(stage_9_per_in[53]),
    .inData_54(stage_9_per_in[54]),
    .inData_55(stage_9_per_in[55]),
    .inData_56(stage_9_per_in[56]),
    .inData_57(stage_9_per_in[57]),
    .inData_58(stage_9_per_in[58]),
    .inData_59(stage_9_per_in[59]),
    .inData_60(stage_9_per_in[60]),
    .inData_61(stage_9_per_in[61]),
    .inData_62(stage_9_per_in[62]),
    .inData_63(stage_9_per_in[63]),
    .outData_0(stage_9_per_out[0]),
    .outData_1(stage_9_per_out[1]),
    .outData_2(stage_9_per_out[2]),
    .outData_3(stage_9_per_out[3]),
    .outData_4(stage_9_per_out[4]),
    .outData_5(stage_9_per_out[5]),
    .outData_6(stage_9_per_out[6]),
    .outData_7(stage_9_per_out[7]),
    .outData_8(stage_9_per_out[8]),
    .outData_9(stage_9_per_out[9]),
    .outData_10(stage_9_per_out[10]),
    .outData_11(stage_9_per_out[11]),
    .outData_12(stage_9_per_out[12]),
    .outData_13(stage_9_per_out[13]),
    .outData_14(stage_9_per_out[14]),
    .outData_15(stage_9_per_out[15]),
    .outData_16(stage_9_per_out[16]),
    .outData_17(stage_9_per_out[17]),
    .outData_18(stage_9_per_out[18]),
    .outData_19(stage_9_per_out[19]),
    .outData_20(stage_9_per_out[20]),
    .outData_21(stage_9_per_out[21]),
    .outData_22(stage_9_per_out[22]),
    .outData_23(stage_9_per_out[23]),
    .outData_24(stage_9_per_out[24]),
    .outData_25(stage_9_per_out[25]),
    .outData_26(stage_9_per_out[26]),
    .outData_27(stage_9_per_out[27]),
    .outData_28(stage_9_per_out[28]),
    .outData_29(stage_9_per_out[29]),
    .outData_30(stage_9_per_out[30]),
    .outData_31(stage_9_per_out[31]),
    .outData_32(stage_9_per_out[32]),
    .outData_33(stage_9_per_out[33]),
    .outData_34(stage_9_per_out[34]),
    .outData_35(stage_9_per_out[35]),
    .outData_36(stage_9_per_out[36]),
    .outData_37(stage_9_per_out[37]),
    .outData_38(stage_9_per_out[38]),
    .outData_39(stage_9_per_out[39]),
    .outData_40(stage_9_per_out[40]),
    .outData_41(stage_9_per_out[41]),
    .outData_42(stage_9_per_out[42]),
    .outData_43(stage_9_per_out[43]),
    .outData_44(stage_9_per_out[44]),
    .outData_45(stage_9_per_out[45]),
    .outData_46(stage_9_per_out[46]),
    .outData_47(stage_9_per_out[47]),
    .outData_48(stage_9_per_out[48]),
    .outData_49(stage_9_per_out[49]),
    .outData_50(stage_9_per_out[50]),
    .outData_51(stage_9_per_out[51]),
    .outData_52(stage_9_per_out[52]),
    .outData_53(stage_9_per_out[53]),
    .outData_54(stage_9_per_out[54]),
    .outData_55(stage_9_per_out[55]),
    .outData_56(stage_9_per_out[56]),
    .outData_57(stage_9_per_out[57]),
    .outData_58(stage_9_per_out[58]),
    .outData_59(stage_9_per_out[59]),
    .outData_60(stage_9_per_out[60]),
    .outData_61(stage_9_per_out[61]),
    .outData_62(stage_9_per_out[62]),
    .outData_63(stage_9_per_out[63]),
    .in_start(in_start[9]),
    .out_start(out_start[9]),
    .clk(clk),
    .rst(rst)
  );

  // TODO(Tian): stage 9 32 butterfly units
  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_0 (
    .x_in(stage_9_per_out[0]),
    .y_in(stage_9_per_out[1]),
    .x_out(outData[0]),
    .y_out(outData[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_1 (
    .x_in(stage_9_per_out[2]),
    .y_in(stage_9_per_out[3]),
    .x_out(outData[2]),
    .y_out(outData[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_2 (
    .x_in(stage_9_per_out[4]),
    .y_in(stage_9_per_out[5]),
    .x_out(outData[4]),
    .y_out(outData[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_3 (
    .x_in(stage_9_per_out[6]),
    .y_in(stage_9_per_out[7]),
    .x_out(outData[6]),
    .y_out(outData[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_4 (
    .x_in(stage_9_per_out[8]),
    .y_in(stage_9_per_out[9]),
    .x_out(outData[8]),
    .y_out(outData[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_5 (
    .x_in(stage_9_per_out[10]),
    .y_in(stage_9_per_out[11]),
    .x_out(outData[10]),
    .y_out(outData[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_6 (
    .x_in(stage_9_per_out[12]),
    .y_in(stage_9_per_out[13]),
    .x_out(outData[12]),
    .y_out(outData[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_7 (
    .x_in(stage_9_per_out[14]),
    .y_in(stage_9_per_out[15]),
    .x_out(outData[14]),
    .y_out(outData[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_8 (
    .x_in(stage_9_per_out[16]),
    .y_in(stage_9_per_out[17]),
    .x_out(outData[16]),
    .y_out(outData[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_9 (
    .x_in(stage_9_per_out[18]),
    .y_in(stage_9_per_out[19]),
    .x_out(outData[18]),
    .y_out(outData[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_10 (
    .x_in(stage_9_per_out[20]),
    .y_in(stage_9_per_out[21]),
    .x_out(outData[20]),
    .y_out(outData[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_11 (
    .x_in(stage_9_per_out[22]),
    .y_in(stage_9_per_out[23]),
    .x_out(outData[22]),
    .y_out(outData[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_12 (
    .x_in(stage_9_per_out[24]),
    .y_in(stage_9_per_out[25]),
    .x_out(outData[24]),
    .y_out(outData[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_13 (
    .x_in(stage_9_per_out[26]),
    .y_in(stage_9_per_out[27]),
    .x_out(outData[26]),
    .y_out(outData[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_14 (
    .x_in(stage_9_per_out[28]),
    .y_in(stage_9_per_out[29]),
    .x_out(outData[28]),
    .y_out(outData[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_15 (
    .x_in(stage_9_per_out[30]),
    .y_in(stage_9_per_out[31]),
    .x_out(outData[30]),
    .y_out(outData[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_16 (
    .x_in(stage_9_per_out[32]),
    .y_in(stage_9_per_out[33]),
    .x_out(outData[32]),
    .y_out(outData[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_17 (
    .x_in(stage_9_per_out[34]),
    .y_in(stage_9_per_out[35]),
    .x_out(outData[34]),
    .y_out(outData[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_18 (
    .x_in(stage_9_per_out[36]),
    .y_in(stage_9_per_out[37]),
    .x_out(outData[36]),
    .y_out(outData[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_19 (
    .x_in(stage_9_per_out[38]),
    .y_in(stage_9_per_out[39]),
    .x_out(outData[38]),
    .y_out(outData[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_20 (
    .x_in(stage_9_per_out[40]),
    .y_in(stage_9_per_out[41]),
    .x_out(outData[40]),
    .y_out(outData[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_21 (
    .x_in(stage_9_per_out[42]),
    .y_in(stage_9_per_out[43]),
    .x_out(outData[42]),
    .y_out(outData[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_22 (
    .x_in(stage_9_per_out[44]),
    .y_in(stage_9_per_out[45]),
    .x_out(outData[44]),
    .y_out(outData[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_23 (
    .x_in(stage_9_per_out[46]),
    .y_in(stage_9_per_out[47]),
    .x_out(outData[46]),
    .y_out(outData[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_24 (
    .x_in(stage_9_per_out[48]),
    .y_in(stage_9_per_out[49]),
    .x_out(outData[48]),
    .y_out(outData[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_25 (
    .x_in(stage_9_per_out[50]),
    .y_in(stage_9_per_out[51]),
    .x_out(outData[50]),
    .y_out(outData[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_26 (
    .x_in(stage_9_per_out[52]),
    .y_in(stage_9_per_out[53]),
    .x_out(outData[52]),
    .y_out(outData[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_27 (
    .x_in(stage_9_per_out[54]),
    .y_in(stage_9_per_out[55]),
    .x_out(outData[54]),
    .y_out(outData[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_28 (
    .x_in(stage_9_per_out[56]),
    .y_in(stage_9_per_out[57]),
    .x_out(outData[56]),
    .y_out(outData[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_29 (
    .x_in(stage_9_per_out[58]),
    .y_in(stage_9_per_out[59]),
    .x_out(outData[58]),
    .y_out(outData[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_30 (
    .x_in(stage_9_per_out[60]),
    .y_in(stage_9_per_out[61]),
    .x_out(outData[60]),
    .y_out(outData[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_31 (
    .x_in(stage_9_per_out[62]),
    .y_in(stage_9_per_out[63]),
    .x_out(outData[62]),
    .y_out(outData[63]),
    .clk(clk),
    .rst(rst)
  );

endmodule
