// NTT Accelerator

module NTT_Top #(
    parameter DATA_WIDTH_PER_INPUT = 28,
    parameter INPUT_PER_CYCLE = 128
  ) (
    inData,
    outData,
    in_start,
    out_start,
    clk,
    rst,
  );

  input clk, rst;

  input in_start[10:0];
  output logic out_start[10:0];

  input        [DATA_WIDTH_PER_INPUT-1:0] inData[INPUT_PER_CYCLE-1:0];
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_0_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_0_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_1_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_1_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_2_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_2_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_3_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_3_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_4_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_4_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_5_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_5_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_6_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_6_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_7_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_7_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_8_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_8_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_9_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_9_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_10_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_10_per_out[INPUT_PER_CYCLE-1:0];

  parameter [7:0] START_CYCLE[12] = {0, 7, 14, 21, 28, 35, 42, 67, 93, 121, 153, 193};

  // TODO(Tian): stage 0 32 butterfly units
  butterfly #(
    .start(START_CYCLE[0]),
    .factors({62736, 248258143, 141200910, 210432655, 60410137, 60657405, 120438379, 154088507,
              168799557, 163194978, 90751938, 174394830, 65612009, 26268761, 42684255, 178512370,
              8259075, 229881708, 81393489, 184579826, 66137976, 168246811, 131575231, 114248229,
              104041706, 39123511, 110271140, 151231163, 9497918, 10785136, 146990305, 228578092}))
  stage_0_butterfly_0 (
    .x_in(inData[0]),
    .y_in(inData[1]),
    .x_out(stage_0_per_in[0]),
    .y_out(stage_0_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({1907454, 179300118, 190023698, 238852009, 90459251, 188631715, 93000404, 68711843,
              145932355, 136072729, 125408694, 234613484, 18646649, 241285957, 249490832, 138558999,
              224650429, 75771663, 118813697, 184231755, 48524018, 184001594, 149996455, 9255299,
              70352813, 49444600, 34248663, 236243144, 125590824, 135108737, 176139969, 129357001}))
  stage_0_butterfly_1 (
    .x_in(inData[2]),
    .y_in(inData[3]),
    .x_out(stage_0_per_in[2]),
    .y_out(stage_0_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({127608977, 157389868, 238966374, 172782070, 127870778, 249304086, 229943365, 896607,
              111929529, 41726718, 264371342, 198700251, 140808004, 155953488, 105651651, 95350060,
              190509603, 169809008, 251686044, 218474935, 65316150, 179814135, 122737973, 239606434,
              221042295, 186854087, 15301013, 24230656, 104126955, 72034061, 83950689, 184896958}))
  stage_0_butterfly_2 (
    .x_in(inData[4]),
    .y_in(inData[5]),
    .x_out(stage_0_per_in[4]),
    .y_out(stage_0_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({169184935, 195652857, 91778054, 32605484, 129584651, 223960411, 35630094, 255719214,
              123658638, 202025824, 210012123, 140340588, 170942291, 215941659, 132315280, 102742547,
              180416915, 30247571, 104447750, 197344625, 194219704, 32737194, 188122907, 179717207,
              72945707, 210644544, 249388588, 181705475, 107928332, 77051365, 46671057, 12667818}))
  stage_0_butterfly_3 (
    .x_in(inData[6]),
    .y_in(inData[7]),
    .x_out(stage_0_per_in[6]),
    .y_out(stage_0_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({221849129, 74962493, 40496733, 229751485, 173052617, 254027033, 200934478, 77856633,
              41023501, 61497280, 230823778, 170978026, 132556999, 24970434, 136104512, 61680409,
              143100858, 163860332, 181610634, 76430728, 181981633, 98483239, 207033531, 228091235,
              8255313, 200339141, 170921357, 158126817, 38773847, 171975768, 247783732, 69921988}))
  stage_0_butterfly_4 (
    .x_in(inData[8]),
    .y_in(inData[9]),
    .x_out(stage_0_per_in[8]),
    .y_out(stage_0_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({172988180, 67529023, 41146808, 88521257, 90342181, 203523838, 234989972, 49058740,
              51002920, 18305869, 67916891, 225077819, 72252210, 143573525, 81013691, 243451530,
              124282928, 198223, 18803294, 253464518, 129798040, 185094855, 265171130, 160882583,
              62374498, 154596247, 168351315, 263412265, 118482368, 248278309, 26045295, 36987199}))
  stage_0_butterfly_5 (
    .x_in(inData[10]),
    .y_in(inData[11]),
    .x_out(stage_0_per_in[10]),
    .y_out(stage_0_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({163149532, 144055138, 120515996, 55158081, 69936597, 215111514, 44459414, 150205042,
              227615757, 246680455, 6265971, 110327668, 50475029, 259992880, 65760618, 161245819,
              87220148, 39654333, 81207363, 7447708, 81762412, 120134099, 252263799, 71887650,
              122977291, 519479, 59384117, 118024210, 110162160, 79702710, 17550542, 132702632}))
  stage_0_butterfly_6 (
    .x_in(inData[12]),
    .y_in(inData[13]),
    .x_out(stage_0_per_in[12]),
    .y_out(stage_0_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({196855462, 205246482, 131370540, 68756958, 97670877, 39872790, 162528302, 170882254,
              138161289, 200939178, 234685655, 210089549, 258291717, 105582618, 176214933, 57174663,
              7092568, 37710032, 267102876, 145439741, 162088178, 193601964, 37647978, 221029739,
              7571096, 23520122, 225275209, 164281505, 156290837, 1058331, 173307030, 100165037}))
  stage_0_butterfly_7 (
    .x_in(inData[14]),
    .y_in(inData[15]),
    .x_out(stage_0_per_in[14]),
    .y_out(stage_0_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({58836748, 229152485, 37016200, 30197592, 198671577, 155288254, 75750547, 151080366,
              24825033, 244557461, 164519211, 98922830, 53079368, 244197291, 144216104, 189539329,
              215423485, 99315902, 196350608, 206880652, 187622314, 15282852, 191761352, 57198083,
              228922625, 245682235, 149687609, 135933105, 90978272, 14827383, 264868967, 222406475}))
  stage_0_butterfly_8 (
    .x_in(inData[16]),
    .y_in(inData[17]),
    .x_out(stage_0_per_in[16]),
    .y_out(stage_0_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({214715735, 196177971, 240473245, 180175431, 238901161, 199052238, 56018142, 99860276,
              142361011, 182231238, 223844182, 250127237, 231138525, 247510253, 150440065, 158154241,
              71354371, 151814684, 14667453, 243146642, 58468223, 94554508, 250276575, 215943874,
              158081289, 101905032, 51995938, 82860468, 264370556, 235758123, 103662145, 183106668}))
  stage_0_butterfly_9 (
    .x_in(inData[18]),
    .y_in(inData[19]),
    .x_out(stage_0_per_in[18]),
    .y_out(stage_0_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({102340758, 129084525, 183756330, 57131388, 39614141, 256641060, 36695937, 74424009,
              173921335, 233895150, 237799186, 252406953, 21531862, 40943954, 20254495, 21576501,
              164861991, 70654895, 101813716, 152512971, 42011142, 166506519, 251811489, 25877458,
              181180691, 94423638, 147769827, 115791483, 242430855, 164243806, 124253615, 157152581}))
  stage_0_butterfly_10 (
    .x_in(inData[20]),
    .y_in(inData[21]),
    .x_out(stage_0_per_in[20]),
    .y_out(stage_0_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({143786732, 149881682, 107655283, 81142751, 159482341, 134571988, 110693156, 185341670,
              15577361, 180088236, 183904649, 195538071, 256986339, 255534095, 45130170, 129933587,
              88993292, 30549918, 39931217, 88157673, 259337446, 51111850, 256691758, 107087275,
              231263484, 264251329, 103488513, 172857441, 11569899, 164573784, 158386056, 65110284}))
  stage_0_butterfly_11 (
    .x_in(inData[22]),
    .y_in(inData[23]),
    .x_out(stage_0_per_in[22]),
    .y_out(stage_0_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({98227373, 29023980, 161075491, 23882789, 22558678, 122229583, 74718485, 104073065,
              128356119, 38864951, 178784227, 173580392, 207607705, 119226838, 155144532, 208507211,
              239045807, 154170583, 84715346, 2673613, 214985679, 113130535, 22397447, 201302943,
              220005950, 241396543, 174624298, 77968856, 68807490, 209917670, 217428510, 193565392}))
  stage_0_butterfly_12 (
    .x_in(inData[24]),
    .y_in(inData[25]),
    .x_out(stage_0_per_in[24]),
    .y_out(stage_0_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({150057464, 23448732, 101070463, 63098068, 209153008, 144072998, 247373572, 210239547,
              122550241, 183262830, 71749872, 180231688, 134429657, 42021864, 12808954, 128052742,
              126302082, 6014167, 78210348, 252922274, 182834104, 201087126, 31027015, 42785182,
              33967221, 48087349, 181325168, 139454911, 212592244, 170346650, 108779799, 89733363}))
  stage_0_butterfly_13 (
    .x_in(inData[26]),
    .y_in(inData[27]),
    .x_out(stage_0_per_in[26]),
    .y_out(stage_0_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({39962754, 256558777, 229530055, 76671502, 260875356, 10696564, 25642441, 109410131,
              53554883, 103692636, 116165973, 51440403, 266139878, 216328989, 173030765, 114527376,
              184347612, 32820960, 176100532, 165433235, 163077087, 89278624, 256453055, 149191288,
              197994960, 138451058, 138996529, 151037716, 49876629, 220416699, 1235353, 183088464}))
  stage_0_butterfly_14 (
    .x_in(inData[28]),
    .y_in(inData[29]),
    .x_out(stage_0_per_in[28]),
    .y_out(stage_0_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({93261610, 172289773, 254832984, 258988459, 108081889, 255307412, 240106988, 231600531,
              159792872, 94389433, 126904432, 211721600, 53728083, 91288416, 78692480, 122077322,
              16344528, 88484653, 187760701, 132336250, 203097121, 158896498, 185758640, 215878737,
              39817818, 36500136, 34527937, 116889475, 138868638, 196733737, 251183310, 167274958}))
  stage_0_butterfly_15 (
    .x_in(inData[30]),
    .y_in(inData[31]),
    .x_out(stage_0_per_in[30]),
    .y_out(stage_0_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({138390585, 237695631, 260020495, 47407140, 50557363, 63634221, 126074738, 131255494,
              209093018, 214996992, 159528330, 39518152, 221285249, 71341164, 171732518, 73723002,
              69789389, 114463563, 219691960, 262334367, 229237307, 253577157, 127322073, 126370638,
              103557733, 187113601, 55682893, 256536575, 123998976, 258162508, 228964332, 108727234}))
  stage_0_butterfly_16 (
    .x_in(inData[32]),
    .y_in(inData[33]),
    .x_out(stage_0_per_in[32]),
    .y_out(stage_0_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({18568532, 142538555, 73697328, 53030863, 148940015, 148753884, 35553140, 249640388,
              196709411, 252862876, 194605816, 241597278, 121142478, 206826789, 147507351, 240078055,
              229741385, 196341244, 217792655, 120846747, 86285917, 182145624, 48555419, 2353936,
              160793918, 110273227, 126498799, 136554164, 57499821, 53524475, 86892569, 244434992}))
  stage_0_butterfly_17 (
    .x_in(inData[34]),
    .y_in(inData[35]),
    .x_out(stage_0_per_in[34]),
    .y_out(stage_0_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({5473511, 144769477, 46912433, 26866408, 213245383, 85422012, 150130406, 169515998,
              132349487, 221059178, 11959677, 219029055, 9479322, 27115908, 36246851, 212385093,
              130771778, 163019788, 107104549, 107135677, 44515532, 263884483, 162829016, 251425486,
              87325743, 211366667, 86460683, 151221429, 11703135, 106563970, 177264548, 225116841}))
  stage_0_butterfly_18 (
    .x_in(inData[36]),
    .y_in(inData[37]),
    .x_out(stage_0_per_in[36]),
    .y_out(stage_0_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({125480909, 5231854, 81083779, 265950738, 81873483, 4986407, 155163691, 208653574,
              112142792, 96892627, 55192006, 60603436, 155517338, 260087354, 90006293, 242826313,
              100132307, 210363951, 164529221, 202640881, 256480283, 123317306, 6725515, 218852619,
              135171113, 9249520, 128889378, 242671835, 48777982, 30822536, 188656071, 56125789}))
  stage_0_butterfly_19 (
    .x_in(inData[38]),
    .y_in(inData[39]),
    .x_out(stage_0_per_in[38]),
    .y_out(stage_0_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({234869713, 226595737, 206537906, 189986560, 42053510, 211444110, 208159538, 242184182,
              234287689, 76639397, 228971558, 245369685, 41652472, 95816060, 82875459, 259733399,
              186545936, 261016176, 243862110, 112718220, 50106798, 84901432, 229222177, 90105969,
              266284483, 148796874, 135646873, 148098547, 166068773, 244602309, 99177320, 255918779}))
  stage_0_butterfly_20 (
    .x_in(inData[40]),
    .y_in(inData[41]),
    .x_out(stage_0_per_in[40]),
    .y_out(stage_0_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({250606181, 149138685, 240784947, 158533760, 212167090, 228871862, 205287356, 61691447,
              109505067, 35559942, 240649845, 62782868, 159471860, 235388028, 230143339, 143816111,
              12651571, 244905743, 175334429, 59370938, 58677377, 249212399, 225914175, 38752877,
              236327891, 157430256, 233906629, 20877990, 220394580, 198378776, 265616179, 260374016}))
  stage_0_butterfly_21 (
    .x_in(inData[42]),
    .y_in(inData[43]),
    .x_out(stage_0_per_in[42]),
    .y_out(stage_0_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({5740730, 218879515, 116970950, 104949331, 42733910, 197423642, 128505750, 96976591,
              151704879, 154775650, 109376139, 162925843, 31551002, 13842453, 181725973, 132907662,
              63656435, 230967163, 149477651, 185120393, 234954565, 46729148, 24734017, 108647642,
              150283834, 67046513, 136400329, 28935497, 99410963, 134843781, 108704486, 41112252}))
  stage_0_butterfly_22 (
    .x_in(inData[44]),
    .y_in(inData[45]),
    .x_out(stage_0_per_in[44]),
    .y_out(stage_0_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({179625763, 21458183, 88419162, 81930, 70436067, 184608754, 39140268, 211152508,
              234322267, 111908324, 243297654, 78892295, 246940389, 192516565, 194815301, 147106083,
              88702124, 59212137, 159725962, 145355888, 35430665, 27694231, 180249606, 70151518,
              21742303, 212770879, 106511467, 171241703, 231268416, 187415781, 138920976, 179287997}))
  stage_0_butterfly_23 (
    .x_in(inData[46]),
    .y_in(inData[47]),
    .x_out(stage_0_per_in[46]),
    .y_out(stage_0_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({106056773, 208950205, 239404299, 263982663, 240039943, 57437223, 100943177, 4470762,
              136599943, 18792168, 179831843, 212470099, 7369182, 144151142, 116861206, 134997518,
              50402804, 45294283, 124269051, 168938760, 159543175, 25904197, 223537938, 151696189,
              106146355, 213752765, 3104477, 204917473, 152734723, 89201641, 10598408, 164702238}))
  stage_0_butterfly_24 (
    .x_in(inData[48]),
    .y_in(inData[49]),
    .x_out(stage_0_per_in[48]),
    .y_out(stage_0_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({58136368, 201838233, 170979076, 63162591, 83840449, 248573392, 225546029, 15349425,
              177927774, 201356021, 113458040, 6044206, 184067420, 70489814, 136415646, 204076371,
              118651137, 98566622, 125694138, 107070533, 250060684, 90061976, 47826324, 226717406,
              61116726, 120964758, 136046821, 165567634, 169435715, 24603905, 123887389, 55517835}))
  stage_0_butterfly_25 (
    .x_in(inData[50]),
    .y_in(inData[51]),
    .x_out(stage_0_per_in[50]),
    .y_out(stage_0_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({104423755, 189611269, 21594518, 225369254, 264479828, 16955107, 183488163, 179315380,
              27503451, 171672871, 122367942, 104310584, 33019077, 156153949, 241508336, 205242093,
              195906424, 9245191, 184151583, 236547476, 67287217, 129666909, 172140914, 176366269,
              188909348, 230339059, 16063721, 54766528, 241821884, 254310437, 210853880, 221585216}))
  stage_0_butterfly_26 (
    .x_in(inData[52]),
    .y_in(inData[53]),
    .x_out(stage_0_per_in[52]),
    .y_out(stage_0_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({136664320, 224508026, 92366490, 78969227, 139852785, 204252016, 106354792, 168672066,
              81860583, 111274912, 133008104, 99112512, 99821278, 34336755, 216240230, 69177824,
              181033780, 59669292, 245310720, 138198441, 106129670, 101060936, 105408561, 129184142,
              194876189, 74816213, 71660202, 185723977, 205958875, 83294274, 242290819, 163860385}))
  stage_0_butterfly_27 (
    .x_in(inData[54]),
    .y_in(inData[55]),
    .x_out(stage_0_per_in[54]),
    .y_out(stage_0_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({63355713, 224551623, 89303497, 59001681, 265709143, 58605619, 6291440, 146899744,
              260400385, 209546662, 184276602, 234070704, 102903513, 224670583, 45907501, 56939589,
              65941195, 93988508, 68363059, 19830371, 85558096, 141580746, 98503463, 160170338,
              79129285, 124727876, 291007, 255492938, 237882452, 8009648, 127215407, 83000954}))
  stage_0_butterfly_28 (
    .x_in(inData[56]),
    .y_in(inData[57]),
    .x_out(stage_0_per_in[56]),
    .y_out(stage_0_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({101375441, 83959851, 142276463, 228944741, 147276523, 175168807, 22914950, 137992276,
              130985550, 198284911, 175012394, 152315952, 118213444, 4622329, 153503748, 225486456,
              107657151, 216371534, 136530068, 35417568, 105733032, 7430278, 41771488, 30147565,
              258487225, 32948426, 177554441, 68094050, 149425076, 117454680, 82939526, 117458270}))
  stage_0_butterfly_29 (
    .x_in(inData[58]),
    .y_in(inData[59]),
    .x_out(stage_0_per_in[58]),
    .y_out(stage_0_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({173776705, 130521421, 149796825, 167654012, 69963660, 242086614, 154162735, 163943008,
              96784305, 178609958, 183166375, 264712232, 42583023, 237453043, 68847542, 245228415,
              17252496, 20606850, 97520605, 151289170, 111517965, 41328094, 140190159, 82596723,
              268107376, 92713113, 217198560, 44239577, 163847221, 13484173, 48025256, 95081716}))
  stage_0_butterfly_30 (
    .x_in(inData[60]),
    .y_in(inData[61]),
    .x_out(stage_0_per_in[60]),
    .y_out(stage_0_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({99627052, 36284828, 193094875, 106508361, 178085825, 67348921, 120761900, 247160596,
              150225643, 241625831, 139998882, 267141235, 249903585, 259081121, 134859556, 163361339,
              26620819, 32461064, 98179318, 213289884, 226850270, 68554215, 216246538, 124135460,
              74278900, 97283065, 118163582, 159360601, 192889387, 65815578, 58580381, 239548624}))
  stage_0_butterfly_31 (
    .x_in(inData[62]),
    .y_in(inData[63]),
    .x_out(stage_0_per_in[62]),
    .y_out(stage_0_per_in[63]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({229351752, 5986200, 238271990, 139336311, 227274721, 217306794, 125625707, 162143577,
              115574858, 4369826, 24738255, 21511271, 151945076, 224561048, 135812431, 96512966,
              86907964, 233570711, 136863777, 193086087, 46407972, 9971642, 215932086, 132028761,
              228870065, 173212060, 130565708, 147718178, 131123953, 167082925, 12430538, 263121861}))
  stage_0_butterfly_32 (
    .x_in(inData[64]),
    .y_in(inData[65]),
    .x_out(stage_0_per_in[64]),
    .y_out(stage_0_per_in[65]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({18284087, 3778321, 215835949, 79816727, 38780522, 180949546, 179673158, 48588607,
              25746466, 68336365, 31768873, 42275209, 82056103, 195819103, 22776264, 241947117,
              132709741, 106442355, 213823426, 222306946, 6841080, 59811701, 108455048, 122257237,
              244570986, 48810421, 35295690, 231200794, 182424131, 84704450, 232516826, 17124429}))
  stage_0_butterfly_33 (
    .x_in(inData[66]),
    .y_in(inData[67]),
    .x_out(stage_0_per_in[66]),
    .y_out(stage_0_per_in[67]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({121332251, 3052481, 154495952, 49806007, 70554670, 54418504, 135886727, 41484727,
              235715975, 27836602, 149329993, 228606302, 25249547, 212109347, 24888645, 158561039,
              260134415, 236342274, 130863524, 244025737, 51724689, 47156256, 108348559, 183216854,
              267488469, 198490305, 97252224, 109429555, 7378856, 140793205, 254596309, 27247099}))
  stage_0_butterfly_34 (
    .x_in(inData[68]),
    .y_in(inData[69]),
    .x_out(stage_0_per_in[68]),
    .y_out(stage_0_per_in[69]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({106831467, 14448911, 36311778, 152480704, 110996066, 45577523, 68771072, 48342959,
              154830655, 121686109, 260828874, 245765723, 125238212, 20537000, 129408474, 44845193,
              237936557, 122360079, 5132066, 13810215, 162923321, 103204044, 217085295, 92792804,
              143112792, 152283243, 60682421, 33223660, 119835732, 150857390, 122169973, 34847782}))
  stage_0_butterfly_35 (
    .x_in(inData[70]),
    .y_in(inData[71]),
    .x_out(stage_0_per_in[70]),
    .y_out(stage_0_per_in[71]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({151923798, 133797910, 2862602, 117960054, 105948718, 20059876, 26464113, 182951273,
              34644106, 265346073, 131105010, 44078325, 47307859, 79305722, 205576016, 192247464,
              233222120, 134390440, 153531059, 101462472, 232770856, 57501675, 46461494, 24794247,
              238036964, 59294895, 118725672, 110117913, 167554606, 84361140, 188917923, 78030852}))
  stage_0_butterfly_36 (
    .x_in(inData[72]),
    .y_in(inData[73]),
    .x_out(stage_0_per_in[72]),
    .y_out(stage_0_per_in[73]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({185050869, 104771116, 129899073, 225676034, 243834156, 156432226, 116017893, 247983171,
              255155441, 12986586, 231410375, 215954984, 112561771, 227071465, 119190794, 60134449,
              131237870, 249630983, 201861189, 107586283, 186098576, 239753050, 158309971, 192193505,
              219418748, 32372991, 33508832, 106358666, 157437159, 38642987, 248241093, 144111858}))
  stage_0_butterfly_37 (
    .x_in(inData[74]),
    .y_in(inData[75]),
    .x_out(stage_0_per_in[74]),
    .y_out(stage_0_per_in[75]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({94277220, 228780544, 12984872, 157537739, 63986967, 171719097, 184499901, 152039665,
              110912131, 182209928, 223045283, 235787722, 36214289, 14462331, 54697818, 259993096,
              68196879, 199075664, 76114224, 120912967, 106463701, 227158983, 170302338, 228212013,
              144673958, 123713876, 178886927, 199074208, 112635657, 213908547, 93347053, 17823318}))
  stage_0_butterfly_38 (
    .x_in(inData[76]),
    .y_in(inData[77]),
    .x_out(stage_0_per_in[76]),
    .y_out(stage_0_per_in[77]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({128643267, 224318864, 131972043, 205821112, 34174616, 265191298, 51441041, 171967455,
              3764785, 113870289, 66804322, 218637579, 92763586, 222708254, 234300746, 259999423,
              79425600, 39822794, 242814722, 108148659, 194119116, 28536923, 57720967, 195919352,
              227038693, 28811566, 161625502, 122116963, 185167965, 117333915, 193454786, 83862241}))
  stage_0_butterfly_39 (
    .x_in(inData[78]),
    .y_in(inData[79]),
    .x_out(stage_0_per_in[78]),
    .y_out(stage_0_per_in[79]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({155464901, 255568559, 757759, 130707805, 137536510, 237348335, 141768337, 223003866,
              176371562, 217608608, 183965087, 267382061, 49387461, 64306041, 30614038, 119248989,
              42144250, 221060093, 208391395, 31181321, 169601951, 131574531, 68378584, 146240700,
              209673396, 51270543, 233335722, 49462279, 8257788, 212712674, 239144038, 126093548}))
  stage_0_butterfly_40 (
    .x_in(inData[80]),
    .y_in(inData[81]),
    .x_out(stage_0_per_in[80]),
    .y_out(stage_0_per_in[81]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({235762007, 205271224, 211663060, 109711544, 16804445, 95429977, 174653765, 104275953,
              214327170, 39463122, 260789685, 130842873, 32828004, 60661841, 155312683, 149391390,
              230428614, 106186088, 69502239, 215911494, 262471786, 101824639, 131432446, 225035437,
              192333550, 8718982, 15958207, 71806036, 232696276, 60363770, 262883371, 41823032}))
  stage_0_butterfly_41 (
    .x_in(inData[82]),
    .y_in(inData[83]),
    .x_out(stage_0_per_in[82]),
    .y_out(stage_0_per_in[83]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({160425732, 189138314, 139937724, 157541500, 225441652, 97602587, 190364932, 43784819,
              244546293, 67840088, 164954582, 238836046, 62948694, 110250618, 109921777, 123166625,
              67538787, 152866160, 194581013, 206403026, 250005524, 224168732, 138660240, 14626898,
              135180292, 164438829, 38284008, 195002054, 195655909, 5958674, 192960909, 219422045}))
  stage_0_butterfly_42 (
    .x_in(inData[84]),
    .y_in(inData[85]),
    .x_out(stage_0_per_in[84]),
    .y_out(stage_0_per_in[85]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({75642576, 257328955, 234828316, 174801883, 112432362, 114891230, 122092755, 59653503,
              229528882, 76662541, 159491283, 204649844, 87947919, 6777444, 48856734, 15637687,
              81695275, 261699407, 237626776, 190689455, 16392555, 163665671, 218881712, 72197923,
              243770087, 48869357, 202431138, 99585718, 170722015, 63257907, 152845826, 214283023}))
  stage_0_butterfly_43 (
    .x_in(inData[86]),
    .y_in(inData[87]),
    .x_out(stage_0_per_in[86]),
    .y_out(stage_0_per_in[87]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({26796856, 166961287, 162545174, 26873848, 264550106, 157511077, 246646236, 103787038,
              29220817, 118901157, 13711872, 156914260, 198369788, 240151518, 95898316, 148505031,
              172925747, 97938637, 34838492, 122693765, 61883556, 65736109, 231672458, 110197348,
              32796042, 207300441, 240095534, 89434836, 49704806, 221163181, 117652871, 86822274}))
  stage_0_butterfly_44 (
    .x_in(inData[88]),
    .y_in(inData[89]),
    .x_out(stage_0_per_in[88]),
    .y_out(stage_0_per_in[89]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({192174913, 205181101, 200114, 187534499, 188446087, 77858155, 78932104, 268045200,
              54047719, 86866558, 245038497, 2963416, 113738086, 247726047, 77729422, 212184418,
              108404040, 160990548, 192227833, 162344188, 225219172, 239353906, 127805784, 259103093,
              263029881, 169234006, 23443169, 77508945, 240905155, 51005918, 83563004, 193603540}))
  stage_0_butterfly_45 (
    .x_in(inData[90]),
    .y_in(inData[91]),
    .x_out(stage_0_per_in[90]),
    .y_out(stage_0_per_in[91]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({83421235, 14751178, 110070131, 71449616, 160647513, 217600940, 260649789, 175074447,
              114016424, 213474870, 179512630, 188754097, 51323950, 247259809, 65690883, 222486214,
              116203844, 33884144, 5695672, 140975706, 135684892, 101029591, 106059530, 23651884,
              119415929, 141473040, 26132679, 12259140, 145011041, 148939130, 135766208, 212842425}))
  stage_0_butterfly_46 (
    .x_in(inData[92]),
    .y_in(inData[93]),
    .x_out(stage_0_per_in[92]),
    .y_out(stage_0_per_in[93]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({141812320, 197944250, 27854761, 5510115, 126711917, 59249925, 86311355, 103407625,
              266701659, 212384234, 55935675, 52557249, 205947916, 50951254, 154254400, 56197115,
              81573675, 117319528, 95352696, 21476942, 80678005, 21249308, 258599303, 114109699,
              44100750, 23918814, 258759731, 95430596, 11447146, 103235635, 180375437, 58071796}))
  stage_0_butterfly_47 (
    .x_in(inData[94]),
    .y_in(inData[95]),
    .x_out(stage_0_per_in[94]),
    .y_out(stage_0_per_in[95]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({232397550, 76613625, 251656189, 30182006, 225306517, 173443464, 115237475, 75233812,
              85762236, 59403344, 174916329, 238064453, 16499278, 81430431, 202855239, 2615849,
              1371159, 196480564, 139897823, 199105134, 49661599, 33454619, 360580, 85118780,
              215247918, 172102431, 234938972, 13664359, 18799530, 242453874, 197777956, 261712272}))
  stage_0_butterfly_48 (
    .x_in(inData[96]),
    .y_in(inData[97]),
    .x_out(stage_0_per_in[96]),
    .y_out(stage_0_per_in[97]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({173978412, 183539945, 35857213, 202544817, 152136534, 107281991, 220692949, 135453164,
              145101039, 56280600, 236121751, 254006109, 267007570, 41756449, 87928571, 13493318,
              21489734, 187504892, 247808775, 28244848, 208868555, 79440456, 16609890, 59625292,
              1618864, 205236559, 46583536, 99167958, 74632878, 167937680, 167199557, 142049175}))
  stage_0_butterfly_49 (
    .x_in(inData[98]),
    .y_in(inData[99]),
    .x_out(stage_0_per_in[98]),
    .y_out(stage_0_per_in[99]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({266521776, 21572447, 56987360, 94223513, 20426733, 66819851, 181022773, 203722503,
              75105065, 2011982, 129605716, 7229020, 206462525, 234710989, 107677384, 194562323,
              49717914, 66144131, 173951180, 246477773, 251263130, 185730304, 14692215, 255690434,
              112251860, 158126231, 153141493, 229582731, 100946881, 34699254, 149344309, 151842442}))
  stage_0_butterfly_50 (
    .x_in(inData[100]),
    .y_in(inData[101]),
    .x_out(stage_0_per_in[100]),
    .y_out(stage_0_per_in[101]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({184791819, 151524267, 56333048, 179139190, 186348595, 8297893, 109371065, 213678319,
              174632895, 258549338, 194603131, 28116292, 66449840, 255738903, 188542273, 78592957,
              5068353, 96374025, 29805745, 197497401, 231677557, 230350716, 69230198, 4491002,
              116647317, 244555167, 90584256, 47508483, 179869441, 175007080, 43714082, 136274746}))
  stage_0_butterfly_51 (
    .x_in(inData[102]),
    .y_in(inData[103]),
    .x_out(stage_0_per_in[102]),
    .y_out(stage_0_per_in[103]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({260851907, 42776728, 39521553, 194846985, 15379209, 61891902, 254332699, 192707093,
              105706660, 152738846, 37752789, 142898101, 158858535, 145592959, 185232992, 204313060,
              260923957, 134614101, 176789033, 97251575, 13704349, 222748125, 109746000, 263215622,
              69414413, 42275800, 207530553, 69218942, 53167918, 150154963, 110104975, 57302073}))
  stage_0_butterfly_52 (
    .x_in(inData[104]),
    .y_in(inData[105]),
    .x_out(stage_0_per_in[104]),
    .y_out(stage_0_per_in[105]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({29470818, 54233307, 132129988, 248896168, 27029386, 26659480, 176832880, 258883039,
              21131779, 66715025, 229784592, 115679885, 153682120, 59375296, 186483628, 72475326,
              157068444, 54358169, 260001724, 209246609, 113781795, 77840672, 179365619, 7116217,
              263718984, 158711864, 74385386, 198306293, 152365066, 245615084, 192872385, 72549374}))
  stage_0_butterfly_53 (
    .x_in(inData[106]),
    .y_in(inData[107]),
    .x_out(stage_0_per_in[106]),
    .y_out(stage_0_per_in[107]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({167586303, 112058009, 63216411, 132200486, 83981669, 12855237, 171842488, 96526884,
              27233477, 264329231, 82632268, 21764948, 144184457, 235284227, 83931467, 97581367,
              136382259, 2029098, 254244111, 102116116, 227944808, 89270439, 213642756, 212003953,
              61250374, 2557700, 170944566, 202918045, 206482017, 235546264, 117771098, 220194496}))
  stage_0_butterfly_54 (
    .x_in(inData[108]),
    .y_in(inData[109]),
    .x_out(stage_0_per_in[108]),
    .y_out(stage_0_per_in[109]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({148827249, 1696019, 58280814, 131559431, 192680584, 13429213, 39919904, 115525972,
              213843114, 17233293, 262250139, 173572777, 162490819, 82054424, 108661782, 157468594,
              97492082, 234121810, 156378126, 185671812, 164207528, 78696193, 204398753, 99516991,
              116801865, 230635721, 15750398, 202001175, 130387641, 37225330, 18191490, 159562860}))
  stage_0_butterfly_55 (
    .x_in(inData[110]),
    .y_in(inData[111]),
    .x_out(stage_0_per_in[110]),
    .y_out(stage_0_per_in[111]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({48491280, 6668530, 24825329, 185532067, 136783171, 211688613, 209177739, 41306715,
              24132582, 146607869, 111072250, 208828758, 171197489, 168472713, 58714599, 206941931,
              183351284, 44427932, 233581580, 130959181, 215737735, 84557377, 165004785, 10658994,
              7620297, 223629100, 165252821, 38635824, 264133989, 76772605, 141503129, 166754761}))
  stage_0_butterfly_56 (
    .x_in(inData[112]),
    .y_in(inData[113]),
    .x_out(stage_0_per_in[112]),
    .y_out(stage_0_per_in[113]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({268021045, 155885829, 194935198, 103408097, 216659963, 190439637, 155010430, 239742054,
              66663233, 179809501, 201979579, 206641346, 127364429, 14129846, 53126633, 134053105,
              111920700, 132259857, 231794807, 157805049, 227465231, 27951846, 168435324, 246208472,
              235669313, 52189384, 40354434, 131200140, 203745198, 13532798, 237430063, 23085612}))
  stage_0_butterfly_57 (
    .x_in(inData[114]),
    .y_in(inData[115]),
    .x_out(stage_0_per_in[114]),
    .y_out(stage_0_per_in[115]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({68227492, 73017801, 9880764, 156474406, 127467506, 169350110, 32128041, 60805498,
              52676293, 83253386, 172273878, 223368694, 83749497, 56381879, 138905259, 221722750,
              107691461, 51218933, 137830340, 232729335, 195074984, 4952604, 16462324, 55752506,
              253757449, 73689066, 169231043, 205614247, 95072757, 264371786, 230124651, 207505578}))
  stage_0_butterfly_58 (
    .x_in(inData[116]),
    .y_in(inData[117]),
    .x_out(stage_0_per_in[116]),
    .y_out(stage_0_per_in[117]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({135770551, 92074820, 203810197, 91588944, 62704870, 236052416, 259685293, 171138130,
              134876482, 55730854, 152468473, 26767263, 92092447, 168849030, 87141435, 96021565,
              201880574, 160584715, 2176252, 248617642, 180394230, 229121016, 171482266, 183002860,
              40301047, 73137377, 28921814, 152308098, 30940476, 154688443, 144681042, 234273255}))
  stage_0_butterfly_59 (
    .x_in(inData[118]),
    .y_in(inData[119]),
    .x_out(stage_0_per_in[118]),
    .y_out(stage_0_per_in[119]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({198563101, 244373783, 198839540, 227953669, 135413478, 118174461, 36389566, 213475348,
              245230909, 170534402, 158032303, 190758660, 115048608, 203514552, 62285640, 150485586,
              43314683, 265006255, 197478524, 110482921, 67824335, 135142897, 174146267, 183449518,
              96257044, 218509565, 227652594, 148811231, 74916156, 251093184, 140577689, 34079608}))
  stage_0_butterfly_60 (
    .x_in(inData[120]),
    .y_in(inData[121]),
    .x_out(stage_0_per_in[120]),
    .y_out(stage_0_per_in[121]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({95052731, 112531453, 85927424, 215784466, 167238213, 230885966, 196216182, 19847969,
              249112263, 215285662, 178662179, 154802450, 40802701, 201888697, 113731328, 68532350,
              200590842, 255059903, 214972665, 202258967, 23130727, 246714101, 208345113, 23277706,
              117177606, 57795922, 161226237, 82689315, 195813478, 44226281, 208881897, 171515704}))
  stage_0_butterfly_61 (
    .x_in(inData[122]),
    .y_in(inData[123]),
    .x_out(stage_0_per_in[122]),
    .y_out(stage_0_per_in[123]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({37560959, 218305863, 37761143, 25592978, 177400482, 125945553, 88343680, 41373747,
              27425418, 99694466, 239054686, 137079211, 177007616, 237567768, 200029177, 257632808,
              236356015, 148722321, 50703780, 113484891, 26760307, 11562888, 224658359, 130055322,
              625780, 215495577, 89497967, 211488291, 216947907, 246176063, 42743336, 76694868}))
  stage_0_butterfly_62 (
    .x_in(inData[124]),
    .y_in(inData[125]),
    .x_out(stage_0_per_in[124]),
    .y_out(stage_0_per_in[125]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({17746678, 145182880, 235736575, 228413454, 10710243, 216347827, 45256937, 32751373,
              143680187, 192995301, 168382927, 139421138, 209077448, 103000049, 3595020, 99532395,
              134045502, 83014713, 91252917, 250977019, 17172477, 101673356, 161740894, 90052819,
              17691838, 266251087, 213947035, 134709760, 1741916, 45566469, 107220558, 127926589}))
  stage_0_butterfly_63 (
    .x_in(inData[126]),
    .y_in(inData[127]),
    .x_out(stage_0_per_in[126]),
    .y_out(stage_0_per_in[127]),
    .clk(clk),
    .rst(rst)
  );




  // TODO(Yang): stage 0 -> stage 1 permutation
  // FIXME: ignore butterfly units for now.
  stage_0_permutation #(
    .DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    .INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_0_1_per (
    .inData_0(stage_0_per_in[0]),
    .inData_1(stage_0_per_in[1]),
    .inData_2(stage_0_per_in[2]),
    .inData_3(stage_0_per_in[3]),
    .inData_4(stage_0_per_in[4]),
    .inData_5(stage_0_per_in[5]),
    .inData_6(stage_0_per_in[6]),
    .inData_7(stage_0_per_in[7]),
    .inData_8(stage_0_per_in[8]),
    .inData_9(stage_0_per_in[9]),
    .inData_10(stage_0_per_in[10]),
    .inData_11(stage_0_per_in[11]),
    .inData_12(stage_0_per_in[12]),
    .inData_13(stage_0_per_in[13]),
    .inData_14(stage_0_per_in[14]),
    .inData_15(stage_0_per_in[15]),
    .inData_16(stage_0_per_in[16]),
    .inData_17(stage_0_per_in[17]),
    .inData_18(stage_0_per_in[18]),
    .inData_19(stage_0_per_in[19]),
    .inData_20(stage_0_per_in[20]),
    .inData_21(stage_0_per_in[21]),
    .inData_22(stage_0_per_in[22]),
    .inData_23(stage_0_per_in[23]),
    .inData_24(stage_0_per_in[24]),
    .inData_25(stage_0_per_in[25]),
    .inData_26(stage_0_per_in[26]),
    .inData_27(stage_0_per_in[27]),
    .inData_28(stage_0_per_in[28]),
    .inData_29(stage_0_per_in[29]),
    .inData_30(stage_0_per_in[30]),
    .inData_31(stage_0_per_in[31]),
    .inData_32(stage_0_per_in[32]),
    .inData_33(stage_0_per_in[33]),
    .inData_34(stage_0_per_in[34]),
    .inData_35(stage_0_per_in[35]),
    .inData_36(stage_0_per_in[36]),
    .inData_37(stage_0_per_in[37]),
    .inData_38(stage_0_per_in[38]),
    .inData_39(stage_0_per_in[39]),
    .inData_40(stage_0_per_in[40]),
    .inData_41(stage_0_per_in[41]),
    .inData_42(stage_0_per_in[42]),
    .inData_43(stage_0_per_in[43]),
    .inData_44(stage_0_per_in[44]),
    .inData_45(stage_0_per_in[45]),
    .inData_46(stage_0_per_in[46]),
    .inData_47(stage_0_per_in[47]),
    .inData_48(stage_0_per_in[48]),
    .inData_49(stage_0_per_in[49]),
    .inData_50(stage_0_per_in[50]),
    .inData_51(stage_0_per_in[51]),
    .inData_52(stage_0_per_in[52]),
    .inData_53(stage_0_per_in[53]),
    .inData_54(stage_0_per_in[54]),
    .inData_55(stage_0_per_in[55]),
    .inData_56(stage_0_per_in[56]),
    .inData_57(stage_0_per_in[57]),
    .inData_58(stage_0_per_in[58]),
    .inData_59(stage_0_per_in[59]),
    .inData_60(stage_0_per_in[60]),
    .inData_61(stage_0_per_in[61]),
    .inData_62(stage_0_per_in[62]),
    .inData_63(stage_0_per_in[63]),
    .inData_64(stage_0_per_in[64]),
    .inData_65(stage_0_per_in[65]),
    .inData_66(stage_0_per_in[66]),
    .inData_67(stage_0_per_in[67]),
    .inData_68(stage_0_per_in[68]),
    .inData_69(stage_0_per_in[69]),
    .inData_70(stage_0_per_in[70]),
    .inData_71(stage_0_per_in[71]),
    .inData_72(stage_0_per_in[72]),
    .inData_73(stage_0_per_in[73]),
    .inData_74(stage_0_per_in[74]),
    .inData_75(stage_0_per_in[75]),
    .inData_76(stage_0_per_in[76]),
    .inData_77(stage_0_per_in[77]),
    .inData_78(stage_0_per_in[78]),
    .inData_79(stage_0_per_in[79]),
    .inData_80(stage_0_per_in[80]),
    .inData_81(stage_0_per_in[81]),
    .inData_82(stage_0_per_in[82]),
    .inData_83(stage_0_per_in[83]),
    .inData_84(stage_0_per_in[84]),
    .inData_85(stage_0_per_in[85]),
    .inData_86(stage_0_per_in[86]),
    .inData_87(stage_0_per_in[87]),
    .inData_88(stage_0_per_in[88]),
    .inData_89(stage_0_per_in[89]),
    .inData_90(stage_0_per_in[90]),
    .inData_91(stage_0_per_in[91]),
    .inData_92(stage_0_per_in[92]),
    .inData_93(stage_0_per_in[93]),
    .inData_94(stage_0_per_in[94]),
    .inData_95(stage_0_per_in[95]),
    .inData_96(stage_0_per_in[96]),
    .inData_97(stage_0_per_in[97]),
    .inData_98(stage_0_per_in[98]),
    .inData_99(stage_0_per_in[99]),
    .inData_100(stage_0_per_in[100]),
    .inData_101(stage_0_per_in[101]),
    .inData_102(stage_0_per_in[102]),
    .inData_103(stage_0_per_in[103]),
    .inData_104(stage_0_per_in[104]),
    .inData_105(stage_0_per_in[105]),
    .inData_106(stage_0_per_in[106]),
    .inData_107(stage_0_per_in[107]),
    .inData_108(stage_0_per_in[108]),
    .inData_109(stage_0_per_in[109]),
    .inData_110(stage_0_per_in[110]),
    .inData_111(stage_0_per_in[111]),
    .inData_112(stage_0_per_in[112]),
    .inData_113(stage_0_per_in[113]),
    .inData_114(stage_0_per_in[114]),
    .inData_115(stage_0_per_in[115]),
    .inData_116(stage_0_per_in[116]),
    .inData_117(stage_0_per_in[117]),
    .inData_118(stage_0_per_in[118]),
    .inData_119(stage_0_per_in[119]),
    .inData_120(stage_0_per_in[120]),
    .inData_121(stage_0_per_in[121]),
    .inData_122(stage_0_per_in[122]),
    .inData_123(stage_0_per_in[123]),
    .inData_124(stage_0_per_in[124]),
    .inData_125(stage_0_per_in[125]),
    .inData_126(stage_0_per_in[126]),
    .inData_127(stage_0_per_in[127]),
    .outData_0(stage_0_per_out[0]),
    .outData_1(stage_0_per_out[1]),
    .outData_2(stage_0_per_out[2]),
    .outData_3(stage_0_per_out[3]),
    .outData_4(stage_0_per_out[4]),
    .outData_5(stage_0_per_out[5]),
    .outData_6(stage_0_per_out[6]),
    .outData_7(stage_0_per_out[7]),
    .outData_8(stage_0_per_out[8]),
    .outData_9(stage_0_per_out[9]),
    .outData_10(stage_0_per_out[10]),
    .outData_11(stage_0_per_out[11]),
    .outData_12(stage_0_per_out[12]),
    .outData_13(stage_0_per_out[13]),
    .outData_14(stage_0_per_out[14]),
    .outData_15(stage_0_per_out[15]),
    .outData_16(stage_0_per_out[16]),
    .outData_17(stage_0_per_out[17]),
    .outData_18(stage_0_per_out[18]),
    .outData_19(stage_0_per_out[19]),
    .outData_20(stage_0_per_out[20]),
    .outData_21(stage_0_per_out[21]),
    .outData_22(stage_0_per_out[22]),
    .outData_23(stage_0_per_out[23]),
    .outData_24(stage_0_per_out[24]),
    .outData_25(stage_0_per_out[25]),
    .outData_26(stage_0_per_out[26]),
    .outData_27(stage_0_per_out[27]),
    .outData_28(stage_0_per_out[28]),
    .outData_29(stage_0_per_out[29]),
    .outData_30(stage_0_per_out[30]),
    .outData_31(stage_0_per_out[31]),
    .outData_32(stage_0_per_out[32]),
    .outData_33(stage_0_per_out[33]),
    .outData_34(stage_0_per_out[34]),
    .outData_35(stage_0_per_out[35]),
    .outData_36(stage_0_per_out[36]),
    .outData_37(stage_0_per_out[37]),
    .outData_38(stage_0_per_out[38]),
    .outData_39(stage_0_per_out[39]),
    .outData_40(stage_0_per_out[40]),
    .outData_41(stage_0_per_out[41]),
    .outData_42(stage_0_per_out[42]),
    .outData_43(stage_0_per_out[43]),
    .outData_44(stage_0_per_out[44]),
    .outData_45(stage_0_per_out[45]),
    .outData_46(stage_0_per_out[46]),
    .outData_47(stage_0_per_out[47]),
    .outData_48(stage_0_per_out[48]),
    .outData_49(stage_0_per_out[49]),
    .outData_50(stage_0_per_out[50]),
    .outData_51(stage_0_per_out[51]),
    .outData_52(stage_0_per_out[52]),
    .outData_53(stage_0_per_out[53]),
    .outData_54(stage_0_per_out[54]),
    .outData_55(stage_0_per_out[55]),
    .outData_56(stage_0_per_out[56]),
    .outData_57(stage_0_per_out[57]),
    .outData_58(stage_0_per_out[58]),
    .outData_59(stage_0_per_out[59]),
    .outData_60(stage_0_per_out[60]),
    .outData_61(stage_0_per_out[61]),
    .outData_62(stage_0_per_out[62]),
    .outData_63(stage_0_per_out[63]),
    .outData_64(stage_0_per_out[64]),
    .outData_65(stage_0_per_out[65]),
    .outData_66(stage_0_per_out[66]),
    .outData_67(stage_0_per_out[67]),
    .outData_68(stage_0_per_out[68]),
    .outData_69(stage_0_per_out[69]),
    .outData_70(stage_0_per_out[70]),
    .outData_71(stage_0_per_out[71]),
    .outData_72(stage_0_per_out[72]),
    .outData_73(stage_0_per_out[73]),
    .outData_74(stage_0_per_out[74]),
    .outData_75(stage_0_per_out[75]),
    .outData_76(stage_0_per_out[76]),
    .outData_77(stage_0_per_out[77]),
    .outData_78(stage_0_per_out[78]),
    .outData_79(stage_0_per_out[79]),
    .outData_80(stage_0_per_out[80]),
    .outData_81(stage_0_per_out[81]),
    .outData_82(stage_0_per_out[82]),
    .outData_83(stage_0_per_out[83]),
    .outData_84(stage_0_per_out[84]),
    .outData_85(stage_0_per_out[85]),
    .outData_86(stage_0_per_out[86]),
    .outData_87(stage_0_per_out[87]),
    .outData_88(stage_0_per_out[88]),
    .outData_89(stage_0_per_out[89]),
    .outData_90(stage_0_per_out[90]),
    .outData_91(stage_0_per_out[91]),
    .outData_92(stage_0_per_out[92]),
    .outData_93(stage_0_per_out[93]),
    .outData_94(stage_0_per_out[94]),
    .outData_95(stage_0_per_out[95]),
    .outData_96(stage_0_per_out[96]),
    .outData_97(stage_0_per_out[97]),
    .outData_98(stage_0_per_out[98]),
    .outData_99(stage_0_per_out[99]),
    .outData_100(stage_0_per_out[100]),
    .outData_101(stage_0_per_out[101]),
    .outData_102(stage_0_per_out[102]),
    .outData_103(stage_0_per_out[103]),
    .outData_104(stage_0_per_out[104]),
    .outData_105(stage_0_per_out[105]),
    .outData_106(stage_0_per_out[106]),
    .outData_107(stage_0_per_out[107]),
    .outData_108(stage_0_per_out[108]),
    .outData_109(stage_0_per_out[109]),
    .outData_110(stage_0_per_out[110]),
    .outData_111(stage_0_per_out[111]),
    .outData_112(stage_0_per_out[112]),
    .outData_113(stage_0_per_out[113]),
    .outData_114(stage_0_per_out[114]),
    .outData_115(stage_0_per_out[115]),
    .outData_116(stage_0_per_out[116]),
    .outData_117(stage_0_per_out[117]),
    .outData_118(stage_0_per_out[118]),
    .outData_119(stage_0_per_out[119]),
    .outData_120(stage_0_per_out[120]),
    .outData_121(stage_0_per_out[121]),
    .outData_122(stage_0_per_out[122]),
    .outData_123(stage_0_per_out[123]),
    .outData_124(stage_0_per_out[124]),
    .outData_125(stage_0_per_out[125]),
    .outData_126(stage_0_per_out[126]),
    .outData_127(stage_0_per_out[127]),
    .in_start(in_start[0]),
    .out_start(out_start[0]),
    .clk(clk),
    .rst(rst)
  );

  // TODO(Tian): stage 1 32 butterfly units
  butterfly #(
    .start(START_CYCLE[1]),
    .factors({178626802, 226568978, 142863934, 100723721, 25937392, 26964940, 49890248, 57740084,
              238700391, 81363847, 185850221, 35411505, 135389110, 34884345, 212020732, 214331009,
              200295213, 154135831, 156023579, 139714595, 214078274, 264282458, 197485473, 167134668,
              245518247, 195063937, 205675156, 251274354, 44349942, 120419308, 75240990, 143647295}))
  stage_1_butterfly_0 (
    .x_in(stage_0_per_out[0]),
    .y_in(stage_0_per_out[1]),
    .x_out(stage_1_per_in[0]),
    .y_out(stage_1_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({178626802, 226568978, 142863934, 100723721, 25937392, 26964940, 49890248, 57740084,
              238700391, 81363847, 185850221, 35411505, 135389110, 34884345, 212020732, 214331009,
              200295213, 154135831, 156023579, 139714595, 214078274, 264282458, 197485473, 167134668,
              245518247, 195063937, 205675156, 251274354, 44349942, 120419308, 75240990, 143647295}))
  stage_1_butterfly_1 (
    .x_in(stage_0_per_out[2]),
    .y_in(stage_0_per_out[3]),
    .x_out(stage_1_per_in[2]),
    .y_out(stage_1_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({241419299, 57439678, 115334054, 66106013, 66456987, 79732409, 185097589, 136199054,
              101221270, 161494327, 227605745, 3059556, 111262804, 170188367, 148511346, 109286034,
              40738286, 180106398, 79909455, 209076586, 107222748, 136983182, 231584900, 145952502,
              260055946, 268223107, 178774268, 5742112, 186303790, 90238900, 135620074, 59970273}))
  stage_1_butterfly_2 (
    .x_in(stage_0_per_out[4]),
    .y_in(stage_0_per_out[5]),
    .x_out(stage_1_per_in[4]),
    .y_out(stage_1_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({241419299, 57439678, 115334054, 66106013, 66456987, 79732409, 185097589, 136199054,
              101221270, 161494327, 227605745, 3059556, 111262804, 170188367, 148511346, 109286034,
              40738286, 180106398, 79909455, 209076586, 107222748, 136983182, 231584900, 145952502,
              260055946, 268223107, 178774268, 5742112, 186303790, 90238900, 135620074, 59970273}))
  stage_1_butterfly_3 (
    .x_in(stage_0_per_out[6]),
    .y_in(stage_0_per_out[7]),
    .x_out(stage_1_per_in[6]),
    .y_out(stage_1_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({202037642, 124029413, 144625416, 152694343, 113912362, 9977836, 194834330, 267034870,
              255819997, 92670067, 10513337, 65501903, 38583127, 219164507, 160223263, 202709135,
              111948379, 158020658, 87171014, 73987125, 71023991, 109238580, 144486207, 156384032,
              66619308, 136306850, 204183192, 37830528, 230038199, 37832342, 184194991, 85850918}))
  stage_1_butterfly_4 (
    .x_in(stage_0_per_out[8]),
    .y_in(stage_0_per_out[9]),
    .x_out(stage_1_per_in[8]),
    .y_out(stage_1_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({202037642, 124029413, 144625416, 152694343, 113912362, 9977836, 194834330, 267034870,
              255819997, 92670067, 10513337, 65501903, 38583127, 219164507, 160223263, 202709135,
              111948379, 158020658, 87171014, 73987125, 71023991, 109238580, 144486207, 156384032,
              66619308, 136306850, 204183192, 37830528, 230038199, 37832342, 184194991, 85850918}))
  stage_1_butterfly_5 (
    .x_in(stage_0_per_out[10]),
    .y_in(stage_0_per_out[11]),
    .x_out(stage_1_per_in[10]),
    .y_out(stage_1_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({224076531, 176876579, 42559975, 181657279, 179710610, 131815160, 22106362, 251982020,
              161018204, 54856389, 141500462, 138344594, 36505175, 107122996, 183471966, 263768524,
              79007221, 75051406, 254205318, 48961458, 236016875, 41046131, 263500442, 238066757,
              173525016, 146660836, 2306944, 233611200, 249749550, 111544693, 216035935, 86146205}))
  stage_1_butterfly_6 (
    .x_in(stage_0_per_out[12]),
    .y_in(stage_0_per_out[13]),
    .x_out(stage_1_per_in[12]),
    .y_out(stage_1_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({224076531, 176876579, 42559975, 181657279, 179710610, 131815160, 22106362, 251982020,
              161018204, 54856389, 141500462, 138344594, 36505175, 107122996, 183471966, 263768524,
              79007221, 75051406, 254205318, 48961458, 236016875, 41046131, 263500442, 238066757,
              173525016, 146660836, 2306944, 233611200, 249749550, 111544693, 216035935, 86146205}))
  stage_1_butterfly_7 (
    .x_in(stage_0_per_out[14]),
    .y_in(stage_0_per_out[15]),
    .x_out(stage_1_per_in[14]),
    .y_out(stage_1_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({262853884, 202016934, 200835165, 139662643, 213369302, 48721923, 77445892, 41376169,
              260565899, 80939041, 28923545, 89821167, 221852517, 116261862, 81165688, 254651521,
              251186267, 173013758, 7373784, 33406019, 256339290, 2568552, 66687, 14131216,
              117147237, 2885885, 69918547, 13809973, 195258296, 232016200, 224618046, 24281843}))
  stage_1_butterfly_8 (
    .x_in(stage_0_per_out[16]),
    .y_in(stage_0_per_out[17]),
    .x_out(stage_1_per_in[16]),
    .y_out(stage_1_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({262853884, 202016934, 200835165, 139662643, 213369302, 48721923, 77445892, 41376169,
              260565899, 80939041, 28923545, 89821167, 221852517, 116261862, 81165688, 254651521,
              251186267, 173013758, 7373784, 33406019, 256339290, 2568552, 66687, 14131216,
              117147237, 2885885, 69918547, 13809973, 195258296, 232016200, 224618046, 24281843}))
  stage_1_butterfly_9 (
    .x_in(stage_0_per_out[18]),
    .y_in(stage_0_per_out[19]),
    .x_out(stage_1_per_in[18]),
    .y_out(stage_1_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({243595082, 205274966, 13214022, 4628244, 204246510, 27222642, 90803899, 156486669,
              2705617, 94113816, 35769351, 180859208, 234383020, 37907807, 82858612, 67895486,
              212990958, 239438610, 82105625, 223749061, 193207980, 22039584, 198659369, 33154381,
              46680870, 57534183, 197375798, 211651639, 85354678, 230913482, 242981970, 118812967}))
  stage_1_butterfly_10 (
    .x_in(stage_0_per_out[20]),
    .y_in(stage_0_per_out[21]),
    .x_out(stage_1_per_in[20]),
    .y_out(stage_1_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({243595082, 205274966, 13214022, 4628244, 204246510, 27222642, 90803899, 156486669,
              2705617, 94113816, 35769351, 180859208, 234383020, 37907807, 82858612, 67895486,
              212990958, 239438610, 82105625, 223749061, 193207980, 22039584, 198659369, 33154381,
              46680870, 57534183, 197375798, 211651639, 85354678, 230913482, 242981970, 118812967}))
  stage_1_butterfly_11 (
    .x_in(stage_0_per_out[22]),
    .y_in(stage_0_per_out[23]),
    .x_out(stage_1_per_in[22]),
    .y_out(stage_1_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({256992454, 239354922, 86047893, 84463383, 174110644, 116219557, 35608242, 28513237,
              230880884, 9083394, 254464819, 63900610, 37207751, 259466327, 258848760, 225061179,
              7004663, 156508649, 193530415, 173627934, 208392312, 161193348, 256317058, 96851793,
              104721465, 188253439, 194631063, 218464636, 175705236, 144500142, 250268531, 208182039}))
  stage_1_butterfly_12 (
    .x_in(stage_0_per_out[24]),
    .y_in(stage_0_per_out[25]),
    .x_out(stage_1_per_in[24]),
    .y_out(stage_1_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({256992454, 239354922, 86047893, 84463383, 174110644, 116219557, 35608242, 28513237,
              230880884, 9083394, 254464819, 63900610, 37207751, 259466327, 258848760, 225061179,
              7004663, 156508649, 193530415, 173627934, 208392312, 161193348, 256317058, 96851793,
              104721465, 188253439, 194631063, 218464636, 175705236, 144500142, 250268531, 208182039}))
  stage_1_butterfly_13 (
    .x_in(stage_0_per_out[26]),
    .y_in(stage_0_per_out[27]),
    .x_out(stage_1_per_in[26]),
    .y_out(stage_1_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({77239454, 143734200, 222855093, 86334506, 21923530, 186026798, 26776855, 42903438,
              58103200, 239780428, 251689720, 253128696, 197145719, 56848151, 164222678, 79432680,
              143288167, 22021280, 248341796, 27523605, 197016099, 171258656, 262755833, 60493834,
              13327732, 14594411, 193102647, 218565763, 57880935, 202657965, 145663803, 68372869}))
  stage_1_butterfly_14 (
    .x_in(stage_0_per_out[28]),
    .y_in(stage_0_per_out[29]),
    .x_out(stage_1_per_in[28]),
    .y_out(stage_1_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({77239454, 143734200, 222855093, 86334506, 21923530, 186026798, 26776855, 42903438,
              58103200, 239780428, 251689720, 253128696, 197145719, 56848151, 164222678, 79432680,
              143288167, 22021280, 248341796, 27523605, 197016099, 171258656, 262755833, 60493834,
              13327732, 14594411, 193102647, 218565763, 57880935, 202657965, 145663803, 68372869}))
  stage_1_butterfly_15 (
    .x_in(stage_0_per_out[30]),
    .y_in(stage_0_per_out[31]),
    .x_out(stage_1_per_in[30]),
    .y_out(stage_1_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({22329094, 146360154, 70370832, 124927121, 43396787, 37292607, 52859373, 41918325,
              224183590, 129161289, 67400723, 48447796, 260125445, 199208092, 157341419, 246555646,
              72618725, 222840723, 116859647, 184120139, 38429557, 253615348, 236609676, 19066791,
              53251080, 41015351, 64307891, 167135704, 254723792, 147133292, 4884476, 124656108}))
  stage_1_butterfly_16 (
    .x_in(stage_0_per_out[32]),
    .y_in(stage_0_per_out[33]),
    .x_out(stage_1_per_in[32]),
    .y_out(stage_1_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({22329094, 146360154, 70370832, 124927121, 43396787, 37292607, 52859373, 41918325,
              224183590, 129161289, 67400723, 48447796, 260125445, 199208092, 157341419, 246555646,
              72618725, 222840723, 116859647, 184120139, 38429557, 253615348, 236609676, 19066791,
              53251080, 41015351, 64307891, 167135704, 254723792, 147133292, 4884476, 124656108}))
  stage_1_butterfly_17 (
    .x_in(stage_0_per_out[34]),
    .y_in(stage_0_per_out[35]),
    .x_out(stage_1_per_in[34]),
    .y_out(stage_1_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({114906207, 93815079, 244981517, 164849679, 182759226, 218411001, 13136617, 248430418,
              48258409, 86611832, 220409117, 98839404, 50041017, 71466452, 6839312, 70993112,
              77785137, 159555178, 168682489, 45900567, 95745785, 266184237, 124689641, 196076822,
              142932928, 26885190, 187973069, 195777196, 242906033, 258128862, 60114085, 203861878}))
  stage_1_butterfly_18 (
    .x_in(stage_0_per_out[36]),
    .y_in(stage_0_per_out[37]),
    .x_out(stage_1_per_in[36]),
    .y_out(stage_1_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({114906207, 93815079, 244981517, 164849679, 182759226, 218411001, 13136617, 248430418,
              48258409, 86611832, 220409117, 98839404, 50041017, 71466452, 6839312, 70993112,
              77785137, 159555178, 168682489, 45900567, 95745785, 266184237, 124689641, 196076822,
              142932928, 26885190, 187973069, 195777196, 242906033, 258128862, 60114085, 203861878}))
  stage_1_butterfly_19 (
    .x_in(stage_0_per_out[38]),
    .y_in(stage_0_per_out[39]),
    .x_out(stage_1_per_in[38]),
    .y_out(stage_1_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({236173805, 59945410, 184394225, 73580010, 38792404, 216197112, 114462613, 264463333,
              127281316, 212643172, 48499686, 67780496, 79121294, 4519531, 233112987, 118263349,
              12994463, 221333762, 252329804, 205553550, 154194427, 246502592, 103784724, 257122505,
              117082039, 85879269, 91384253, 253166836, 222792306, 19111856, 233855133, 74620568}))
  stage_1_butterfly_20 (
    .x_in(stage_0_per_out[40]),
    .y_in(stage_0_per_out[41]),
    .x_out(stage_1_per_in[40]),
    .y_out(stage_1_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({236173805, 59945410, 184394225, 73580010, 38792404, 216197112, 114462613, 264463333,
              127281316, 212643172, 48499686, 67780496, 79121294, 4519531, 233112987, 118263349,
              12994463, 221333762, 252329804, 205553550, 154194427, 246502592, 103784724, 257122505,
              117082039, 85879269, 91384253, 253166836, 222792306, 19111856, 233855133, 74620568}))
  stage_1_butterfly_21 (
    .x_in(stage_0_per_out[42]),
    .y_in(stage_0_per_out[43]),
    .x_out(stage_1_per_in[42]),
    .y_out(stage_1_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({154634100, 195704814, 100279875, 265093046, 64402402, 22419281, 130965208, 239219986,
              185120175, 258398710, 127264350, 205236983, 105759020, 65162419, 199811874, 3615863,
              126437335, 67459976, 178639438, 43817935, 219155874, 209365645, 87333346, 95592544,
              240329350, 83440545, 109752985, 91771920, 252048491, 23196483, 45533578, 153870377}))
  stage_1_butterfly_22 (
    .x_in(stage_0_per_out[44]),
    .y_in(stage_0_per_out[45]),
    .x_out(stage_1_per_in[44]),
    .y_out(stage_1_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({154634100, 195704814, 100279875, 265093046, 64402402, 22419281, 130965208, 239219986,
              185120175, 258398710, 127264350, 205236983, 105759020, 65162419, 199811874, 3615863,
              126437335, 67459976, 178639438, 43817935, 219155874, 209365645, 87333346, 95592544,
              240329350, 83440545, 109752985, 91771920, 252048491, 23196483, 45533578, 153870377}))
  stage_1_butterfly_23 (
    .x_in(stage_0_per_out[46]),
    .y_in(stage_0_per_out[47]),
    .x_out(stage_1_per_in[46]),
    .y_out(stage_1_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({82346526, 58372872, 226865216, 5284602, 30998042, 182147827, 1381761, 57884406,
              126629575, 14425613, 61366355, 234435452, 189834774, 193726599, 224367752, 260962587,
              110001979, 230614882, 90833651, 41031357, 223156719, 102404987, 93188095, 95943159,
              216344829, 77043356, 76840577, 126638229, 175434645, 228233519, 21699914, 149817301}))
  stage_1_butterfly_24 (
    .x_in(stage_0_per_out[48]),
    .y_in(stage_0_per_out[49]),
    .x_out(stage_1_per_in[48]),
    .y_out(stage_1_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({82346526, 58372872, 226865216, 5284602, 30998042, 182147827, 1381761, 57884406,
              126629575, 14425613, 61366355, 234435452, 189834774, 193726599, 224367752, 260962587,
              110001979, 230614882, 90833651, 41031357, 223156719, 102404987, 93188095, 95943159,
              216344829, 77043356, 76840577, 126638229, 175434645, 228233519, 21699914, 149817301}))
  stage_1_butterfly_25 (
    .x_in(stage_0_per_out[50]),
    .y_in(stage_0_per_out[51]),
    .x_out(stage_1_per_in[50]),
    .y_out(stage_1_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({124972666, 35010964, 144113751, 146661492, 248813222, 209335538, 64059298, 95362545,
              12562435, 121954140, 133033169, 176649880, 200991325, 191064173, 11713205, 24417340,
              50422568, 152117270, 209487240, 140766862, 199654780, 237702991, 53666796, 200880844,
              54194127, 53103748, 85925921, 39159482, 82994670, 151554022, 131606898, 185196127}))
  stage_1_butterfly_26 (
    .x_in(stage_0_per_out[52]),
    .y_in(stage_0_per_out[53]),
    .x_out(stage_1_per_in[52]),
    .y_out(stage_1_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({124972666, 35010964, 144113751, 146661492, 248813222, 209335538, 64059298, 95362545,
              12562435, 121954140, 133033169, 176649880, 200991325, 191064173, 11713205, 24417340,
              50422568, 152117270, 209487240, 140766862, 199654780, 237702991, 53666796, 200880844,
              54194127, 53103748, 85925921, 39159482, 82994670, 151554022, 131606898, 185196127}))
  stage_1_butterfly_27 (
    .x_in(stage_0_per_out[54]),
    .y_in(stage_0_per_out[55]),
    .x_out(stage_1_per_in[54]),
    .y_out(stage_1_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({259902883, 32769539, 253791818, 90415400, 141049304, 201671086, 69255389, 148688834,
              5071752, 18362334, 134836604, 239800333, 94872102, 77506253, 124878920, 163120146,
              96098889, 70871651, 242696977, 95276657, 203277373, 28990836, 16822583, 122635188,
              185121114, 225384963, 148548934, 41573703, 231508432, 94729012, 189935724, 243900215}))
  stage_1_butterfly_28 (
    .x_in(stage_0_per_out[56]),
    .y_in(stage_0_per_out[57]),
    .x_out(stage_1_per_in[56]),
    .y_out(stage_1_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({259902883, 32769539, 253791818, 90415400, 141049304, 201671086, 69255389, 148688834,
              5071752, 18362334, 134836604, 239800333, 94872102, 77506253, 124878920, 163120146,
              96098889, 70871651, 242696977, 95276657, 203277373, 28990836, 16822583, 122635188,
              185121114, 225384963, 148548934, 41573703, 231508432, 94729012, 189935724, 243900215}))
  stage_1_butterfly_29 (
    .x_in(stage_0_per_out[58]),
    .y_in(stage_0_per_out[59]),
    .x_out(stage_1_per_in[58]),
    .y_out(stage_1_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({127717239, 6456449, 172630653, 217483488, 137520333, 139730465, 248206642, 22116392,
              259334239, 13394971, 112174110, 179888950, 16703359, 197641184, 143389876, 74661667,
              75588758, 4184358, 33161823, 107466416, 14369566, 243789725, 133797547, 38723858,
              227177249, 215351473, 55952036, 192111834, 186728485, 153057061, 170437415, 6554463}))
  stage_1_butterfly_30 (
    .x_in(stage_0_per_out[60]),
    .y_in(stage_0_per_out[61]),
    .x_out(stage_1_per_in[60]),
    .y_out(stage_1_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({127717239, 6456449, 172630653, 217483488, 137520333, 139730465, 248206642, 22116392,
              259334239, 13394971, 112174110, 179888950, 16703359, 197641184, 143389876, 74661667,
              75588758, 4184358, 33161823, 107466416, 14369566, 243789725, 133797547, 38723858,
              227177249, 215351473, 55952036, 192111834, 186728485, 153057061, 170437415, 6554463}))
  stage_1_butterfly_31 (
    .x_in(stage_0_per_out[62]),
    .y_in(stage_0_per_out[63]),
    .x_out(stage_1_per_in[62]),
    .y_out(stage_1_per_in[63]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({36426289, 228368554, 98446051, 195462811, 48496256, 236960516, 58870518, 148535761,
              170998790, 54281363, 153913781, 90710559, 26451456, 189299702, 50385541, 46629005,
              6208689, 99461488, 47430573, 143466178, 118216948, 173116375, 9453674, 157049837,
              43737855, 264289232, 54092187, 198072981, 100770703, 224620084, 267404879, 133881133}))
  stage_1_butterfly_32 (
    .x_in(stage_0_per_out[64]),
    .y_in(stage_0_per_out[65]),
    .x_out(stage_1_per_in[64]),
    .y_out(stage_1_per_in[65]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({36426289, 228368554, 98446051, 195462811, 48496256, 236960516, 58870518, 148535761,
              170998790, 54281363, 153913781, 90710559, 26451456, 189299702, 50385541, 46629005,
              6208689, 99461488, 47430573, 143466178, 118216948, 173116375, 9453674, 157049837,
              43737855, 264289232, 54092187, 198072981, 100770703, 224620084, 267404879, 133881133}))
  stage_1_butterfly_33 (
    .x_in(stage_0_per_out[66]),
    .y_in(stage_0_per_out[67]),
    .x_out(stage_1_per_in[66]),
    .y_out(stage_1_per_in[67]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({189966412, 104968162, 213018760, 150529015, 266940341, 61436946, 230680452, 72619804,
              65241583, 129726580, 196403691, 262108538, 39377609, 188624074, 175901771, 124518160,
              39161232, 219432305, 259358426, 145040924, 106026444, 119641299, 118804291, 58085086,
              26707009, 141552463, 68124275, 73785583, 89556414, 211474022, 80152118, 78067214}))
  stage_1_butterfly_34 (
    .x_in(stage_0_per_out[68]),
    .y_in(stage_0_per_out[69]),
    .x_out(stage_1_per_in[68]),
    .y_out(stage_1_per_in[69]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({189966412, 104968162, 213018760, 150529015, 266940341, 61436946, 230680452, 72619804,
              65241583, 129726580, 196403691, 262108538, 39377609, 188624074, 175901771, 124518160,
              39161232, 219432305, 259358426, 145040924, 106026444, 119641299, 118804291, 58085086,
              26707009, 141552463, 68124275, 73785583, 89556414, 211474022, 80152118, 78067214}))
  stage_1_butterfly_35 (
    .x_in(stage_0_per_out[70]),
    .y_in(stage_0_per_out[71]),
    .x_out(stage_1_per_in[70]),
    .y_out(stage_1_per_in[71]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({141057137, 258951073, 83042590, 247893310, 153843002, 203299319, 127868408, 90431622,
              190155959, 25148713, 224762304, 72006316, 138773321, 34739971, 60791061, 154200425,
              248800534, 20654843, 84553412, 89839882, 208367077, 140702439, 198469359, 243002151,
              255369977, 27101256, 215044990, 176150397, 84103703, 109081133, 161356640, 61148806}))
  stage_1_butterfly_36 (
    .x_in(stage_0_per_out[72]),
    .y_in(stage_0_per_out[73]),
    .x_out(stage_1_per_in[72]),
    .y_out(stage_1_per_in[73]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({141057137, 258951073, 83042590, 247893310, 153843002, 203299319, 127868408, 90431622,
              190155959, 25148713, 224762304, 72006316, 138773321, 34739971, 60791061, 154200425,
              248800534, 20654843, 84553412, 89839882, 208367077, 140702439, 198469359, 243002151,
              255369977, 27101256, 215044990, 176150397, 84103703, 109081133, 161356640, 61148806}))
  stage_1_butterfly_37 (
    .x_in(stage_0_per_out[74]),
    .y_in(stage_0_per_out[75]),
    .x_out(stage_1_per_in[74]),
    .y_out(stage_1_per_in[75]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({75414331, 55709426, 9179161, 95442771, 188476710, 214979600, 127510598, 217412044,
              82911469, 34957318, 176271587, 207338429, 35544064, 89363633, 79351768, 245466834,
              72719897, 104015737, 77136822, 73243528, 16967674, 205950205, 20490089, 176574100,
              215608734, 207179347, 217413665, 76831465, 131659808, 252140774, 201376724, 115561740}))
  stage_1_butterfly_38 (
    .x_in(stage_0_per_out[76]),
    .y_in(stage_0_per_out[77]),
    .x_out(stage_1_per_in[76]),
    .y_out(stage_1_per_in[77]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({75414331, 55709426, 9179161, 95442771, 188476710, 214979600, 127510598, 217412044,
              82911469, 34957318, 176271587, 207338429, 35544064, 89363633, 79351768, 245466834,
              72719897, 104015737, 77136822, 73243528, 16967674, 205950205, 20490089, 176574100,
              215608734, 207179347, 217413665, 76831465, 131659808, 252140774, 201376724, 115561740}))
  stage_1_butterfly_39 (
    .x_in(stage_0_per_out[78]),
    .y_in(stage_0_per_out[79]),
    .x_out(stage_1_per_in[78]),
    .y_out(stage_1_per_in[79]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({204172184, 144194814, 155441062, 209967729, 193915015, 222818810, 151896708, 207289252,
              192679930, 40189829, 169229772, 74346844, 216420108, 150921330, 172134458, 143985240,
              188623776, 192273850, 202075477, 76213351, 259641163, 94417879, 82259521, 226423252,
              259932536, 232035425, 166849602, 217984510, 144316291, 91036891, 18026307, 168335279}))
  stage_1_butterfly_40 (
    .x_in(stage_0_per_out[80]),
    .y_in(stage_0_per_out[81]),
    .x_out(stage_1_per_in[80]),
    .y_out(stage_1_per_in[81]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({204172184, 144194814, 155441062, 209967729, 193915015, 222818810, 151896708, 207289252,
              192679930, 40189829, 169229772, 74346844, 216420108, 150921330, 172134458, 143985240,
              188623776, 192273850, 202075477, 76213351, 259641163, 94417879, 82259521, 226423252,
              259932536, 232035425, 166849602, 217984510, 144316291, 91036891, 18026307, 168335279}))
  stage_1_butterfly_41 (
    .x_in(stage_0_per_out[82]),
    .y_in(stage_0_per_out[83]),
    .x_out(stage_1_per_in[82]),
    .y_out(stage_1_per_in[83]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({114289273, 80852279, 183986337, 255259435, 146691665, 165177241, 253065021, 182882105,
              171586403, 154399218, 177621090, 27789608, 103427147, 180135303, 111988251, 75455626,
              176645554, 244247525, 197737960, 204890405, 258770065, 7487276, 149046252, 33861678,
              64324001, 212068395, 248421583, 262436297, 239135625, 186920055, 119165597, 88850354}))
  stage_1_butterfly_42 (
    .x_in(stage_0_per_out[84]),
    .y_in(stage_0_per_out[85]),
    .x_out(stage_1_per_in[84]),
    .y_out(stage_1_per_in[85]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({114289273, 80852279, 183986337, 255259435, 146691665, 165177241, 253065021, 182882105,
              171586403, 154399218, 177621090, 27789608, 103427147, 180135303, 111988251, 75455626,
              176645554, 244247525, 197737960, 204890405, 258770065, 7487276, 149046252, 33861678,
              64324001, 212068395, 248421583, 262436297, 239135625, 186920055, 119165597, 88850354}))
  stage_1_butterfly_43 (
    .x_in(stage_0_per_out[86]),
    .y_in(stage_0_per_out[87]),
    .x_out(stage_1_per_in[86]),
    .y_out(stage_1_per_in[87]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({266373219, 34279912, 209875154, 121172029, 250769297, 242437879, 181957723, 25651112,
              207436891, 35697312, 29380441, 34535827, 104305160, 22230677, 245673827, 211697180,
              154780521, 76495986, 113066699, 112847505, 139316176, 184571212, 178875242, 247989601,
              155494097, 147907047, 243436973, 177240151, 138028127, 106663692, 110007683, 78372181}))
  stage_1_butterfly_44 (
    .x_in(stage_0_per_out[88]),
    .y_in(stage_0_per_out[89]),
    .x_out(stage_1_per_in[88]),
    .y_out(stage_1_per_in[89]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({266373219, 34279912, 209875154, 121172029, 250769297, 242437879, 181957723, 25651112,
              207436891, 35697312, 29380441, 34535827, 104305160, 22230677, 245673827, 211697180,
              154780521, 76495986, 113066699, 112847505, 139316176, 184571212, 178875242, 247989601,
              155494097, 147907047, 243436973, 177240151, 138028127, 106663692, 110007683, 78372181}))
  stage_1_butterfly_45 (
    .x_in(stage_0_per_out[90]),
    .y_in(stage_0_per_out[91]),
    .x_out(stage_1_per_in[90]),
    .y_out(stage_1_per_in[91]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({148884778, 236741674, 57044952, 126959268, 126650083, 33343400, 40931981, 63912782,
              166350047, 91136142, 110850189, 81924749, 187446019, 255364493, 124441328, 39292866,
              210949816, 117619035, 123481104, 153827860, 250734390, 106713399, 108936038, 152193297,
              130184658, 260941520, 267667077, 162889363, 98151275, 141192231, 142379740, 252921174}))
  stage_1_butterfly_46 (
    .x_in(stage_0_per_out[92]),
    .y_in(stage_0_per_out[93]),
    .x_out(stage_1_per_in[92]),
    .y_out(stage_1_per_in[93]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({148884778, 236741674, 57044952, 126959268, 126650083, 33343400, 40931981, 63912782,
              166350047, 91136142, 110850189, 81924749, 187446019, 255364493, 124441328, 39292866,
              210949816, 117619035, 123481104, 153827860, 250734390, 106713399, 108936038, 152193297,
              130184658, 260941520, 267667077, 162889363, 98151275, 141192231, 142379740, 252921174}))
  stage_1_butterfly_47 (
    .x_in(stage_0_per_out[94]),
    .y_in(stage_0_per_out[95]),
    .x_out(stage_1_per_in[94]),
    .y_out(stage_1_per_in[95]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({150629496, 175887545, 171269635, 236561162, 213843220, 91188581, 108521058, 67911621,
              104486975, 100791881, 247062782, 211284483, 46126435, 222236846, 31157387, 38115064,
              145706676, 106939991, 264758616, 17337072, 195763450, 3677235, 126894636, 66528431,
              179997990, 81431484, 204816575, 91524025, 75117738, 141917139, 254692251, 45684920}))
  stage_1_butterfly_48 (
    .x_in(stage_0_per_out[96]),
    .y_in(stage_0_per_out[97]),
    .x_out(stage_1_per_in[96]),
    .y_out(stage_1_per_in[97]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({150629496, 175887545, 171269635, 236561162, 213843220, 91188581, 108521058, 67911621,
              104486975, 100791881, 247062782, 211284483, 46126435, 222236846, 31157387, 38115064,
              145706676, 106939991, 264758616, 17337072, 195763450, 3677235, 126894636, 66528431,
              179997990, 81431484, 204816575, 91524025, 75117738, 141917139, 254692251, 45684920}))
  stage_1_butterfly_49 (
    .x_in(stage_0_per_out[98]),
    .y_in(stage_0_per_out[99]),
    .x_out(stage_1_per_in[98]),
    .y_out(stage_1_per_in[99]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({95956458, 119248786, 25402945, 253446904, 65939487, 105651679, 86425411, 104273059,
              32326785, 248049881, 60951044, 128923754, 51590619, 81879124, 50250252, 202017141,
              166705511, 176106545, 99151986, 135965343, 196552678, 36678208, 250979164, 242448751,
              232700332, 157159811, 49412866, 24169593, 123556687, 66398989, 79759830, 47380903}))
  stage_1_butterfly_50 (
    .x_in(stage_0_per_out[100]),
    .y_in(stage_0_per_out[101]),
    .x_out(stage_1_per_in[100]),
    .y_out(stage_1_per_in[101]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({95956458, 119248786, 25402945, 253446904, 65939487, 105651679, 86425411, 104273059,
              32326785, 248049881, 60951044, 128923754, 51590619, 81879124, 50250252, 202017141,
              166705511, 176106545, 99151986, 135965343, 196552678, 36678208, 250979164, 242448751,
              232700332, 157159811, 49412866, 24169593, 123556687, 66398989, 79759830, 47380903}))
  stage_1_butterfly_51 (
    .x_in(stage_0_per_out[102]),
    .y_in(stage_0_per_out[103]),
    .x_out(stage_1_per_in[102]),
    .y_out(stage_1_per_in[103]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({218922070, 88068083, 224193580, 38581987, 22320040, 213462715, 232970901, 143364478,
              167753662, 182920379, 145595829, 120068412, 122372515, 126673466, 267701123, 83665434,
              106279827, 261080375, 115935405, 237391515, 153619107, 248921617, 96644160, 54591848,
              205764394, 230500375, 166918201, 58002164, 174707320, 120623833, 215876710, 117068649}))
  stage_1_butterfly_52 (
    .x_in(stage_0_per_out[104]),
    .y_in(stage_0_per_out[105]),
    .x_out(stage_1_per_in[104]),
    .y_out(stage_1_per_in[105]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({218922070, 88068083, 224193580, 38581987, 22320040, 213462715, 232970901, 143364478,
              167753662, 182920379, 145595829, 120068412, 122372515, 126673466, 267701123, 83665434,
              106279827, 261080375, 115935405, 237391515, 153619107, 248921617, 96644160, 54591848,
              205764394, 230500375, 166918201, 58002164, 174707320, 120623833, 215876710, 117068649}))
  stage_1_butterfly_53 (
    .x_in(stage_0_per_out[106]),
    .y_in(stage_0_per_out[107]),
    .x_out(stage_1_per_in[106]),
    .y_out(stage_1_per_in[107]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({158913333, 176734838, 145325214, 11727916, 60782408, 20002868, 104683412, 123982174,
              254862428, 86422302, 95857789, 63759475, 61255010, 220487343, 253117467, 114664154,
              78726832, 175735543, 104494180, 7525756, 238828812, 21397846, 59853183, 80415871,
              243959994, 44095704, 213675734, 83594289, 215932651, 209775390, 129973973, 177655074}))
  stage_1_butterfly_54 (
    .x_in(stage_0_per_out[108]),
    .y_in(stage_0_per_out[109]),
    .x_out(stage_1_per_in[108]),
    .y_out(stage_1_per_in[109]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({158913333, 176734838, 145325214, 11727916, 60782408, 20002868, 104683412, 123982174,
              254862428, 86422302, 95857789, 63759475, 61255010, 220487343, 253117467, 114664154,
              78726832, 175735543, 104494180, 7525756, 238828812, 21397846, 59853183, 80415871,
              243959994, 44095704, 213675734, 83594289, 215932651, 209775390, 129973973, 177655074}))
  stage_1_butterfly_55 (
    .x_in(stage_0_per_out[110]),
    .y_in(stage_0_per_out[111]),
    .x_out(stage_1_per_in[110]),
    .y_out(stage_1_per_in[111]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({125480758, 128081279, 196727396, 133543242, 53716996, 26713518, 171508784, 5028136,
              267892175, 50106553, 14195884, 73917671, 195995970, 181264550, 79252444, 125264465,
              264722248, 232215778, 18807047, 79343207, 205816155, 192939426, 262718787, 15406607,
              116341913, 148816114, 145444168, 258312618, 175360485, 85861280, 158406994, 146642358}))
  stage_1_butterfly_56 (
    .x_in(stage_0_per_out[112]),
    .y_in(stage_0_per_out[113]),
    .x_out(stage_1_per_in[112]),
    .y_out(stage_1_per_in[113]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({125480758, 128081279, 196727396, 133543242, 53716996, 26713518, 171508784, 5028136,
              267892175, 50106553, 14195884, 73917671, 195995970, 181264550, 79252444, 125264465,
              264722248, 232215778, 18807047, 79343207, 205816155, 192939426, 262718787, 15406607,
              116341913, 148816114, 145444168, 258312618, 175360485, 85861280, 158406994, 146642358}))
  stage_1_butterfly_57 (
    .x_in(stage_0_per_out[114]),
    .y_in(stage_0_per_out[115]),
    .x_out(stage_1_per_in[114]),
    .y_out(stage_1_per_in[115]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({59278718, 48487396, 8772869, 34093582, 140980229, 264638858, 187469377, 70333973,
              100306740, 202839194, 178750844, 132216843, 203006324, 226857524, 6515518, 214119665,
              22483780, 52952054, 119598304, 176646986, 27342032, 80711179, 114157546, 184171973,
              104225870, 85943438, 146917464, 239243318, 24889364, 165873702, 71397785, 159375180}))
  stage_1_butterfly_58 (
    .x_in(stage_0_per_out[116]),
    .y_in(stage_0_per_out[117]),
    .x_out(stage_1_per_in[116]),
    .y_out(stage_1_per_in[117]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({59278718, 48487396, 8772869, 34093582, 140980229, 264638858, 187469377, 70333973,
              100306740, 202839194, 178750844, 132216843, 203006324, 226857524, 6515518, 214119665,
              22483780, 52952054, 119598304, 176646986, 27342032, 80711179, 114157546, 184171973,
              104225870, 85943438, 146917464, 239243318, 24889364, 165873702, 71397785, 159375180}))
  stage_1_butterfly_59 (
    .x_in(stage_0_per_out[118]),
    .y_in(stage_0_per_out[119]),
    .x_out(stage_1_per_in[118]),
    .y_out(stage_1_per_in[119]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({64064097, 136417444, 157208225, 182812696, 144089543, 81774581, 256522921, 212200386,
              50115805, 96014882, 223616593, 241368847, 38129962, 221869909, 119697484, 217885801,
              259065776, 41460117, 25013575, 71010071, 62424622, 18485653, 255875272, 155632772,
              134337294, 139206238, 176530780, 127930513, 73886338, 52942312, 75752194, 4980542}))
  stage_1_butterfly_60 (
    .x_in(stage_0_per_out[120]),
    .y_in(stage_0_per_out[121]),
    .x_out(stage_1_per_in[120]),
    .y_out(stage_1_per_in[121]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({64064097, 136417444, 157208225, 182812696, 144089543, 81774581, 256522921, 212200386,
              50115805, 96014882, 223616593, 241368847, 38129962, 221869909, 119697484, 217885801,
              259065776, 41460117, 25013575, 71010071, 62424622, 18485653, 255875272, 155632772,
              134337294, 139206238, 176530780, 127930513, 73886338, 52942312, 75752194, 4980542}))
  stage_1_butterfly_61 (
    .x_in(stage_0_per_out[122]),
    .y_in(stage_0_per_out[123]),
    .x_out(stage_1_per_in[122]),
    .y_out(stage_1_per_in[123]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({135644103, 157158700, 51299486, 254780782, 50213981, 108532653, 34242638, 134518349,
              152505970, 187892585, 254241553, 256890018, 35688570, 153805373, 258225039, 50021352,
              209423491, 179675005, 31515852, 244217621, 27456585, 94477870, 207692352, 12048336,
              48893661, 102888853, 157311612, 116226, 187345691, 106441080, 126420356, 101380813}))
  stage_1_butterfly_62 (
    .x_in(stage_0_per_out[124]),
    .y_in(stage_0_per_out[125]),
    .x_out(stage_1_per_in[124]),
    .y_out(stage_1_per_in[125]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({135644103, 157158700, 51299486, 254780782, 50213981, 108532653, 34242638, 134518349,
              152505970, 187892585, 254241553, 256890018, 35688570, 153805373, 258225039, 50021352,
              209423491, 179675005, 31515852, 244217621, 27456585, 94477870, 207692352, 12048336,
              48893661, 102888853, 157311612, 116226, 187345691, 106441080, 126420356, 101380813}))
  stage_1_butterfly_63 (
    .x_in(stage_0_per_out[126]),
    .y_in(stage_0_per_out[127]),
    .x_out(stage_1_per_in[126]),
    .y_out(stage_1_per_in[127]),
    .clk(clk),
    .rst(rst)
  );


  
  // TODO(Yang): stage 1 -> stage 2 permutation
  // FIXME: ignore butterfly units for now.
  stage_1_permutation #(
    .DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    .INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_1_2_per (
    .inData_0(stage_1_per_in[0]),
    .inData_1(stage_1_per_in[1]),
    .inData_2(stage_1_per_in[2]),
    .inData_3(stage_1_per_in[3]),
    .inData_4(stage_1_per_in[4]),
    .inData_5(stage_1_per_in[5]),
    .inData_6(stage_1_per_in[6]),
    .inData_7(stage_1_per_in[7]),
    .inData_8(stage_1_per_in[8]),
    .inData_9(stage_1_per_in[9]),
    .inData_10(stage_1_per_in[10]),
    .inData_11(stage_1_per_in[11]),
    .inData_12(stage_1_per_in[12]),
    .inData_13(stage_1_per_in[13]),
    .inData_14(stage_1_per_in[14]),
    .inData_15(stage_1_per_in[15]),
    .inData_16(stage_1_per_in[16]),
    .inData_17(stage_1_per_in[17]),
    .inData_18(stage_1_per_in[18]),
    .inData_19(stage_1_per_in[19]),
    .inData_20(stage_1_per_in[20]),
    .inData_21(stage_1_per_in[21]),
    .inData_22(stage_1_per_in[22]),
    .inData_23(stage_1_per_in[23]),
    .inData_24(stage_1_per_in[24]),
    .inData_25(stage_1_per_in[25]),
    .inData_26(stage_1_per_in[26]),
    .inData_27(stage_1_per_in[27]),
    .inData_28(stage_1_per_in[28]),
    .inData_29(stage_1_per_in[29]),
    .inData_30(stage_1_per_in[30]),
    .inData_31(stage_1_per_in[31]),
    .inData_32(stage_1_per_in[32]),
    .inData_33(stage_1_per_in[33]),
    .inData_34(stage_1_per_in[34]),
    .inData_35(stage_1_per_in[35]),
    .inData_36(stage_1_per_in[36]),
    .inData_37(stage_1_per_in[37]),
    .inData_38(stage_1_per_in[38]),
    .inData_39(stage_1_per_in[39]),
    .inData_40(stage_1_per_in[40]),
    .inData_41(stage_1_per_in[41]),
    .inData_42(stage_1_per_in[42]),
    .inData_43(stage_1_per_in[43]),
    .inData_44(stage_1_per_in[44]),
    .inData_45(stage_1_per_in[45]),
    .inData_46(stage_1_per_in[46]),
    .inData_47(stage_1_per_in[47]),
    .inData_48(stage_1_per_in[48]),
    .inData_49(stage_1_per_in[49]),
    .inData_50(stage_1_per_in[50]),
    .inData_51(stage_1_per_in[51]),
    .inData_52(stage_1_per_in[52]),
    .inData_53(stage_1_per_in[53]),
    .inData_54(stage_1_per_in[54]),
    .inData_55(stage_1_per_in[55]),
    .inData_56(stage_1_per_in[56]),
    .inData_57(stage_1_per_in[57]),
    .inData_58(stage_1_per_in[58]),
    .inData_59(stage_1_per_in[59]),
    .inData_60(stage_1_per_in[60]),
    .inData_61(stage_1_per_in[61]),
    .inData_62(stage_1_per_in[62]),
    .inData_63(stage_1_per_in[63]),
    .inData_64(stage_1_per_in[64]),
    .inData_65(stage_1_per_in[65]),
    .inData_66(stage_1_per_in[66]),
    .inData_67(stage_1_per_in[67]),
    .inData_68(stage_1_per_in[68]),
    .inData_69(stage_1_per_in[69]),
    .inData_70(stage_1_per_in[70]),
    .inData_71(stage_1_per_in[71]),
    .inData_72(stage_1_per_in[72]),
    .inData_73(stage_1_per_in[73]),
    .inData_74(stage_1_per_in[74]),
    .inData_75(stage_1_per_in[75]),
    .inData_76(stage_1_per_in[76]),
    .inData_77(stage_1_per_in[77]),
    .inData_78(stage_1_per_in[78]),
    .inData_79(stage_1_per_in[79]),
    .inData_80(stage_1_per_in[80]),
    .inData_81(stage_1_per_in[81]),
    .inData_82(stage_1_per_in[82]),
    .inData_83(stage_1_per_in[83]),
    .inData_84(stage_1_per_in[84]),
    .inData_85(stage_1_per_in[85]),
    .inData_86(stage_1_per_in[86]),
    .inData_87(stage_1_per_in[87]),
    .inData_88(stage_1_per_in[88]),
    .inData_89(stage_1_per_in[89]),
    .inData_90(stage_1_per_in[90]),
    .inData_91(stage_1_per_in[91]),
    .inData_92(stage_1_per_in[92]),
    .inData_93(stage_1_per_in[93]),
    .inData_94(stage_1_per_in[94]),
    .inData_95(stage_1_per_in[95]),
    .inData_96(stage_1_per_in[96]),
    .inData_97(stage_1_per_in[97]),
    .inData_98(stage_1_per_in[98]),
    .inData_99(stage_1_per_in[99]),
    .inData_100(stage_1_per_in[100]),
    .inData_101(stage_1_per_in[101]),
    .inData_102(stage_1_per_in[102]),
    .inData_103(stage_1_per_in[103]),
    .inData_104(stage_1_per_in[104]),
    .inData_105(stage_1_per_in[105]),
    .inData_106(stage_1_per_in[106]),
    .inData_107(stage_1_per_in[107]),
    .inData_108(stage_1_per_in[108]),
    .inData_109(stage_1_per_in[109]),
    .inData_110(stage_1_per_in[110]),
    .inData_111(stage_1_per_in[111]),
    .inData_112(stage_1_per_in[112]),
    .inData_113(stage_1_per_in[113]),
    .inData_114(stage_1_per_in[114]),
    .inData_115(stage_1_per_in[115]),
    .inData_116(stage_1_per_in[116]),
    .inData_117(stage_1_per_in[117]),
    .inData_118(stage_1_per_in[118]),
    .inData_119(stage_1_per_in[119]),
    .inData_120(stage_1_per_in[120]),
    .inData_121(stage_1_per_in[121]),
    .inData_122(stage_1_per_in[122]),
    .inData_123(stage_1_per_in[123]),
    .inData_124(stage_1_per_in[124]),
    .inData_125(stage_1_per_in[125]),
    .inData_126(stage_1_per_in[126]),
    .inData_127(stage_1_per_in[127]),
    .outData_0(stage_1_per_out[0]),
    .outData_1(stage_1_per_out[1]),
    .outData_2(stage_1_per_out[2]),
    .outData_3(stage_1_per_out[3]),
    .outData_4(stage_1_per_out[4]),
    .outData_5(stage_1_per_out[5]),
    .outData_6(stage_1_per_out[6]),
    .outData_7(stage_1_per_out[7]),
    .outData_8(stage_1_per_out[8]),
    .outData_9(stage_1_per_out[9]),
    .outData_10(stage_1_per_out[10]),
    .outData_11(stage_1_per_out[11]),
    .outData_12(stage_1_per_out[12]),
    .outData_13(stage_1_per_out[13]),
    .outData_14(stage_1_per_out[14]),
    .outData_15(stage_1_per_out[15]),
    .outData_16(stage_1_per_out[16]),
    .outData_17(stage_1_per_out[17]),
    .outData_18(stage_1_per_out[18]),
    .outData_19(stage_1_per_out[19]),
    .outData_20(stage_1_per_out[20]),
    .outData_21(stage_1_per_out[21]),
    .outData_22(stage_1_per_out[22]),
    .outData_23(stage_1_per_out[23]),
    .outData_24(stage_1_per_out[24]),
    .outData_25(stage_1_per_out[25]),
    .outData_26(stage_1_per_out[26]),
    .outData_27(stage_1_per_out[27]),
    .outData_28(stage_1_per_out[28]),
    .outData_29(stage_1_per_out[29]),
    .outData_30(stage_1_per_out[30]),
    .outData_31(stage_1_per_out[31]),
    .outData_32(stage_1_per_out[32]),
    .outData_33(stage_1_per_out[33]),
    .outData_34(stage_1_per_out[34]),
    .outData_35(stage_1_per_out[35]),
    .outData_36(stage_1_per_out[36]),
    .outData_37(stage_1_per_out[37]),
    .outData_38(stage_1_per_out[38]),
    .outData_39(stage_1_per_out[39]),
    .outData_40(stage_1_per_out[40]),
    .outData_41(stage_1_per_out[41]),
    .outData_42(stage_1_per_out[42]),
    .outData_43(stage_1_per_out[43]),
    .outData_44(stage_1_per_out[44]),
    .outData_45(stage_1_per_out[45]),
    .outData_46(stage_1_per_out[46]),
    .outData_47(stage_1_per_out[47]),
    .outData_48(stage_1_per_out[48]),
    .outData_49(stage_1_per_out[49]),
    .outData_50(stage_1_per_out[50]),
    .outData_51(stage_1_per_out[51]),
    .outData_52(stage_1_per_out[52]),
    .outData_53(stage_1_per_out[53]),
    .outData_54(stage_1_per_out[54]),
    .outData_55(stage_1_per_out[55]),
    .outData_56(stage_1_per_out[56]),
    .outData_57(stage_1_per_out[57]),
    .outData_58(stage_1_per_out[58]),
    .outData_59(stage_1_per_out[59]),
    .outData_60(stage_1_per_out[60]),
    .outData_61(stage_1_per_out[61]),
    .outData_62(stage_1_per_out[62]),
    .outData_63(stage_1_per_out[63]),
    .outData_64(stage_1_per_out[64]),
    .outData_65(stage_1_per_out[65]),
    .outData_66(stage_1_per_out[66]),
    .outData_67(stage_1_per_out[67]),
    .outData_68(stage_1_per_out[68]),
    .outData_69(stage_1_per_out[69]),
    .outData_70(stage_1_per_out[70]),
    .outData_71(stage_1_per_out[71]),
    .outData_72(stage_1_per_out[72]),
    .outData_73(stage_1_per_out[73]),
    .outData_74(stage_1_per_out[74]),
    .outData_75(stage_1_per_out[75]),
    .outData_76(stage_1_per_out[76]),
    .outData_77(stage_1_per_out[77]),
    .outData_78(stage_1_per_out[78]),
    .outData_79(stage_1_per_out[79]),
    .outData_80(stage_1_per_out[80]),
    .outData_81(stage_1_per_out[81]),
    .outData_82(stage_1_per_out[82]),
    .outData_83(stage_1_per_out[83]),
    .outData_84(stage_1_per_out[84]),
    .outData_85(stage_1_per_out[85]),
    .outData_86(stage_1_per_out[86]),
    .outData_87(stage_1_per_out[87]),
    .outData_88(stage_1_per_out[88]),
    .outData_89(stage_1_per_out[89]),
    .outData_90(stage_1_per_out[90]),
    .outData_91(stage_1_per_out[91]),
    .outData_92(stage_1_per_out[92]),
    .outData_93(stage_1_per_out[93]),
    .outData_94(stage_1_per_out[94]),
    .outData_95(stage_1_per_out[95]),
    .outData_96(stage_1_per_out[96]),
    .outData_97(stage_1_per_out[97]),
    .outData_98(stage_1_per_out[98]),
    .outData_99(stage_1_per_out[99]),
    .outData_100(stage_1_per_out[100]),
    .outData_101(stage_1_per_out[101]),
    .outData_102(stage_1_per_out[102]),
    .outData_103(stage_1_per_out[103]),
    .outData_104(stage_1_per_out[104]),
    .outData_105(stage_1_per_out[105]),
    .outData_106(stage_1_per_out[106]),
    .outData_107(stage_1_per_out[107]),
    .outData_108(stage_1_per_out[108]),
    .outData_109(stage_1_per_out[109]),
    .outData_110(stage_1_per_out[110]),
    .outData_111(stage_1_per_out[111]),
    .outData_112(stage_1_per_out[112]),
    .outData_113(stage_1_per_out[113]),
    .outData_114(stage_1_per_out[114]),
    .outData_115(stage_1_per_out[115]),
    .outData_116(stage_1_per_out[116]),
    .outData_117(stage_1_per_out[117]),
    .outData_118(stage_1_per_out[118]),
    .outData_119(stage_1_per_out[119]),
    .outData_120(stage_1_per_out[120]),
    .outData_121(stage_1_per_out[121]),
    .outData_122(stage_1_per_out[122]),
    .outData_123(stage_1_per_out[123]),
    .outData_124(stage_1_per_out[124]),
    .outData_125(stage_1_per_out[125]),
    .outData_126(stage_1_per_out[126]),
    .outData_127(stage_1_per_out[127]),
    .in_start(in_start[1]),
    .out_start(out_start[1]),
    .clk(clk),
    .rst(rst)
  );


  // TODO(Tian): stage 2 32 butterfly units
  butterfly #(
    .start(START_CYCLE[2]),
    .factors({187381670, 120217110, 54714468, 142656304, 196018390, 212112171, 26068775, 174191574,
              27439037, 189139684, 58661398, 128297265, 174612628, 23442787, 35629855, 50083600,
              233083676, 24365404, 173628384, 63661975, 142941966, 252714435, 10646661, 156195364,
              250031819, 183613005, 206844979, 78273516, 121414397, 72509307, 255478273, 255463943}))
  stage_2_butterfly_0 (
    .x_in(stage_1_per_out[0]),
    .y_in(stage_1_per_out[1]),
    .x_out(stage_2_per_in[0]),
    .y_out(stage_2_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({187381670, 120217110, 54714468, 142656304, 196018390, 212112171, 26068775, 174191574,
              27439037, 189139684, 58661398, 128297265, 174612628, 23442787, 35629855, 50083600,
              233083676, 24365404, 173628384, 63661975, 142941966, 252714435, 10646661, 156195364,
              250031819, 183613005, 206844979, 78273516, 121414397, 72509307, 255478273, 255463943}))
  stage_2_butterfly_1 (
    .x_in(stage_1_per_out[2]),
    .y_in(stage_1_per_out[3]),
    .x_out(stage_2_per_in[2]),
    .y_out(stage_2_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({187381670, 120217110, 54714468, 142656304, 196018390, 212112171, 26068775, 174191574,
              27439037, 189139684, 58661398, 128297265, 174612628, 23442787, 35629855, 50083600,
              233083676, 24365404, 173628384, 63661975, 142941966, 252714435, 10646661, 156195364,
              250031819, 183613005, 206844979, 78273516, 121414397, 72509307, 255478273, 255463943}))
  stage_2_butterfly_2 (
    .x_in(stage_1_per_out[4]),
    .y_in(stage_1_per_out[5]),
    .x_out(stage_2_per_in[4]),
    .y_out(stage_2_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({187381670, 120217110, 54714468, 142656304, 196018390, 212112171, 26068775, 174191574,
              27439037, 189139684, 58661398, 128297265, 174612628, 23442787, 35629855, 50083600,
              233083676, 24365404, 173628384, 63661975, 142941966, 252714435, 10646661, 156195364,
              250031819, 183613005, 206844979, 78273516, 121414397, 72509307, 255478273, 255463943}))
  stage_2_butterfly_3 (
    .x_in(stage_1_per_out[6]),
    .y_in(stage_1_per_out[7]),
    .x_out(stage_2_per_in[6]),
    .y_out(stage_2_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({222912429, 248922055, 38252193, 157839041, 243009216, 21649526, 187208958, 116527240,
              189909138, 190586128, 224322272, 130154791, 75993973, 259621463, 509728, 190565686,
              82779345, 211982342, 58491201, 147903734, 128589211, 165001005, 267008435, 147014646,
              54690936, 174163034, 53284215, 226025718, 156298941, 73072346, 186048173, 112360014}))
  stage_2_butterfly_4 (
    .x_in(stage_1_per_out[8]),
    .y_in(stage_1_per_out[9]),
    .x_out(stage_2_per_in[8]),
    .y_out(stage_2_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({222912429, 248922055, 38252193, 157839041, 243009216, 21649526, 187208958, 116527240,
              189909138, 190586128, 224322272, 130154791, 75993973, 259621463, 509728, 190565686,
              82779345, 211982342, 58491201, 147903734, 128589211, 165001005, 267008435, 147014646,
              54690936, 174163034, 53284215, 226025718, 156298941, 73072346, 186048173, 112360014}))
  stage_2_butterfly_5 (
    .x_in(stage_1_per_out[10]),
    .y_in(stage_1_per_out[11]),
    .x_out(stage_2_per_in[10]),
    .y_out(stage_2_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({222912429, 248922055, 38252193, 157839041, 243009216, 21649526, 187208958, 116527240,
              189909138, 190586128, 224322272, 130154791, 75993973, 259621463, 509728, 190565686,
              82779345, 211982342, 58491201, 147903734, 128589211, 165001005, 267008435, 147014646,
              54690936, 174163034, 53284215, 226025718, 156298941, 73072346, 186048173, 112360014}))
  stage_2_butterfly_6 (
    .x_in(stage_1_per_out[12]),
    .y_in(stage_1_per_out[13]),
    .x_out(stage_2_per_in[12]),
    .y_out(stage_2_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({222912429, 248922055, 38252193, 157839041, 243009216, 21649526, 187208958, 116527240,
              189909138, 190586128, 224322272, 130154791, 75993973, 259621463, 509728, 190565686,
              82779345, 211982342, 58491201, 147903734, 128589211, 165001005, 267008435, 147014646,
              54690936, 174163034, 53284215, 226025718, 156298941, 73072346, 186048173, 112360014}))
  stage_2_butterfly_7 (
    .x_in(stage_1_per_out[14]),
    .y_in(stage_1_per_out[15]),
    .x_out(stage_2_per_in[14]),
    .y_out(stage_2_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({224391994, 29779638, 217763430, 107830842, 193911793, 168470500, 267506256, 82483914,
              231354349, 133273987, 149788353, 6760936, 54916848, 207530748, 36492987, 91458750,
              202032572, 69017626, 139374293, 268043824, 158314046, 121608761, 153237233, 159491687,
              19700796, 8474832, 81838336, 148491526, 13228372, 255552842, 8836114, 256519333}))
  stage_2_butterfly_8 (
    .x_in(stage_1_per_out[16]),
    .y_in(stage_1_per_out[17]),
    .x_out(stage_2_per_in[16]),
    .y_out(stage_2_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({224391994, 29779638, 217763430, 107830842, 193911793, 168470500, 267506256, 82483914,
              231354349, 133273987, 149788353, 6760936, 54916848, 207530748, 36492987, 91458750,
              202032572, 69017626, 139374293, 268043824, 158314046, 121608761, 153237233, 159491687,
              19700796, 8474832, 81838336, 148491526, 13228372, 255552842, 8836114, 256519333}))
  stage_2_butterfly_9 (
    .x_in(stage_1_per_out[18]),
    .y_in(stage_1_per_out[19]),
    .x_out(stage_2_per_in[18]),
    .y_out(stage_2_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({224391994, 29779638, 217763430, 107830842, 193911793, 168470500, 267506256, 82483914,
              231354349, 133273987, 149788353, 6760936, 54916848, 207530748, 36492987, 91458750,
              202032572, 69017626, 139374293, 268043824, 158314046, 121608761, 153237233, 159491687,
              19700796, 8474832, 81838336, 148491526, 13228372, 255552842, 8836114, 256519333}))
  stage_2_butterfly_10 (
    .x_in(stage_1_per_out[20]),
    .y_in(stage_1_per_out[21]),
    .x_out(stage_2_per_in[20]),
    .y_out(stage_2_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({224391994, 29779638, 217763430, 107830842, 193911793, 168470500, 267506256, 82483914,
              231354349, 133273987, 149788353, 6760936, 54916848, 207530748, 36492987, 91458750,
              202032572, 69017626, 139374293, 268043824, 158314046, 121608761, 153237233, 159491687,
              19700796, 8474832, 81838336, 148491526, 13228372, 255552842, 8836114, 256519333}))
  stage_2_butterfly_11 (
    .x_in(stage_1_per_out[22]),
    .y_in(stage_1_per_out[23]),
    .x_out(stage_2_per_in[22]),
    .y_out(stage_2_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({134161265, 165671105, 184464011, 218207344, 236272786, 33594840, 197065781, 14882191,
              114052864, 129677075, 189757297, 159978713, 171198428, 195152646, 99543252, 94436408,
              36196902, 160050812, 20655050, 145034434, 233967292, 134796549, 184560259, 99012968,
              243047656, 54393228, 94686133, 195270185, 249947221, 132747224, 237395333, 227454343}))
  stage_2_butterfly_12 (
    .x_in(stage_1_per_out[24]),
    .y_in(stage_1_per_out[25]),
    .x_out(stage_2_per_in[24]),
    .y_out(stage_2_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({134161265, 165671105, 184464011, 218207344, 236272786, 33594840, 197065781, 14882191,
              114052864, 129677075, 189757297, 159978713, 171198428, 195152646, 99543252, 94436408,
              36196902, 160050812, 20655050, 145034434, 233967292, 134796549, 184560259, 99012968,
              243047656, 54393228, 94686133, 195270185, 249947221, 132747224, 237395333, 227454343}))
  stage_2_butterfly_13 (
    .x_in(stage_1_per_out[26]),
    .y_in(stage_1_per_out[27]),
    .x_out(stage_2_per_in[26]),
    .y_out(stage_2_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({134161265, 165671105, 184464011, 218207344, 236272786, 33594840, 197065781, 14882191,
              114052864, 129677075, 189757297, 159978713, 171198428, 195152646, 99543252, 94436408,
              36196902, 160050812, 20655050, 145034434, 233967292, 134796549, 184560259, 99012968,
              243047656, 54393228, 94686133, 195270185, 249947221, 132747224, 237395333, 227454343}))
  stage_2_butterfly_14 (
    .x_in(stage_1_per_out[28]),
    .y_in(stage_1_per_out[29]),
    .x_out(stage_2_per_in[28]),
    .y_out(stage_2_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({134161265, 165671105, 184464011, 218207344, 236272786, 33594840, 197065781, 14882191,
              114052864, 129677075, 189757297, 159978713, 171198428, 195152646, 99543252, 94436408,
              36196902, 160050812, 20655050, 145034434, 233967292, 134796549, 184560259, 99012968,
              243047656, 54393228, 94686133, 195270185, 249947221, 132747224, 237395333, 227454343}))
  stage_2_butterfly_15 (
    .x_in(stage_1_per_out[30]),
    .y_in(stage_1_per_out[31]),
    .x_out(stage_2_per_in[30]),
    .y_out(stage_2_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({64830196, 70325928, 163197321, 102034957, 31964447, 251717800, 9205704, 85566308,
              148108490, 237616434, 128052734, 113049121, 261143222, 211201491, 151857114, 53025186,
              74918627, 83194655, 31540722, 167181901, 32160642, 38415865, 264974639, 36213609,
              156534179, 148649408, 42575603, 263102666, 47531240, 212425161, 19817676, 25652741}))
  stage_2_butterfly_16 (
    .x_in(stage_1_per_out[32]),
    .y_in(stage_1_per_out[33]),
    .x_out(stage_2_per_in[32]),
    .y_out(stage_2_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({64830196, 70325928, 163197321, 102034957, 31964447, 251717800, 9205704, 85566308,
              148108490, 237616434, 128052734, 113049121, 261143222, 211201491, 151857114, 53025186,
              74918627, 83194655, 31540722, 167181901, 32160642, 38415865, 264974639, 36213609,
              156534179, 148649408, 42575603, 263102666, 47531240, 212425161, 19817676, 25652741}))
  stage_2_butterfly_17 (
    .x_in(stage_1_per_out[34]),
    .y_in(stage_1_per_out[35]),
    .x_out(stage_2_per_in[34]),
    .y_out(stage_2_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({64830196, 70325928, 163197321, 102034957, 31964447, 251717800, 9205704, 85566308,
              148108490, 237616434, 128052734, 113049121, 261143222, 211201491, 151857114, 53025186,
              74918627, 83194655, 31540722, 167181901, 32160642, 38415865, 264974639, 36213609,
              156534179, 148649408, 42575603, 263102666, 47531240, 212425161, 19817676, 25652741}))
  stage_2_butterfly_18 (
    .x_in(stage_1_per_out[36]),
    .y_in(stage_1_per_out[37]),
    .x_out(stage_2_per_in[36]),
    .y_out(stage_2_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({64830196, 70325928, 163197321, 102034957, 31964447, 251717800, 9205704, 85566308,
              148108490, 237616434, 128052734, 113049121, 261143222, 211201491, 151857114, 53025186,
              74918627, 83194655, 31540722, 167181901, 32160642, 38415865, 264974639, 36213609,
              156534179, 148649408, 42575603, 263102666, 47531240, 212425161, 19817676, 25652741}))
  stage_2_butterfly_19 (
    .x_in(stage_1_per_out[38]),
    .y_in(stage_1_per_out[39]),
    .x_out(stage_2_per_in[38]),
    .y_out(stage_2_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({62456195, 139101859, 18205961, 107513427, 90701762, 228715598, 122609533, 37504237,
              157649589, 102785717, 123720956, 212728405, 163812077, 257402730, 29537138, 248946430,
              129694458, 222087036, 183590673, 111532362, 12711531, 162575967, 86752434, 153316076,
              61348732, 67784869, 168674209, 199055975, 5368199, 37377133, 127918992, 143811089}))
  stage_2_butterfly_20 (
    .x_in(stage_1_per_out[40]),
    .y_in(stage_1_per_out[41]),
    .x_out(stage_2_per_in[40]),
    .y_out(stage_2_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({62456195, 139101859, 18205961, 107513427, 90701762, 228715598, 122609533, 37504237,
              157649589, 102785717, 123720956, 212728405, 163812077, 257402730, 29537138, 248946430,
              129694458, 222087036, 183590673, 111532362, 12711531, 162575967, 86752434, 153316076,
              61348732, 67784869, 168674209, 199055975, 5368199, 37377133, 127918992, 143811089}))
  stage_2_butterfly_21 (
    .x_in(stage_1_per_out[42]),
    .y_in(stage_1_per_out[43]),
    .x_out(stage_2_per_in[42]),
    .y_out(stage_2_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({62456195, 139101859, 18205961, 107513427, 90701762, 228715598, 122609533, 37504237,
              157649589, 102785717, 123720956, 212728405, 163812077, 257402730, 29537138, 248946430,
              129694458, 222087036, 183590673, 111532362, 12711531, 162575967, 86752434, 153316076,
              61348732, 67784869, 168674209, 199055975, 5368199, 37377133, 127918992, 143811089}))
  stage_2_butterfly_22 (
    .x_in(stage_1_per_out[44]),
    .y_in(stage_1_per_out[45]),
    .x_out(stage_2_per_in[44]),
    .y_out(stage_2_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({62456195, 139101859, 18205961, 107513427, 90701762, 228715598, 122609533, 37504237,
              157649589, 102785717, 123720956, 212728405, 163812077, 257402730, 29537138, 248946430,
              129694458, 222087036, 183590673, 111532362, 12711531, 162575967, 86752434, 153316076,
              61348732, 67784869, 168674209, 199055975, 5368199, 37377133, 127918992, 143811089}))
  stage_2_butterfly_23 (
    .x_in(stage_1_per_out[46]),
    .y_in(stage_1_per_out[47]),
    .x_out(stage_2_per_in[46]),
    .y_out(stage_2_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({48885659, 205681680, 46120362, 175949223, 233437339, 127163336, 79843127, 90149574,
              158914825, 248133554, 264322432, 229032903, 7376627, 4643973, 120080647, 98269185,
              92379159, 160048836, 184522009, 254234203, 100343421, 195181845, 66412546, 126749676,
              247452694, 266777211, 12551837, 161345834, 255457916, 59214954, 110302060, 135080569}))
  stage_2_butterfly_24 (
    .x_in(stage_1_per_out[48]),
    .y_in(stage_1_per_out[49]),
    .x_out(stage_2_per_in[48]),
    .y_out(stage_2_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({48885659, 205681680, 46120362, 175949223, 233437339, 127163336, 79843127, 90149574,
              158914825, 248133554, 264322432, 229032903, 7376627, 4643973, 120080647, 98269185,
              92379159, 160048836, 184522009, 254234203, 100343421, 195181845, 66412546, 126749676,
              247452694, 266777211, 12551837, 161345834, 255457916, 59214954, 110302060, 135080569}))
  stage_2_butterfly_25 (
    .x_in(stage_1_per_out[50]),
    .y_in(stage_1_per_out[51]),
    .x_out(stage_2_per_in[50]),
    .y_out(stage_2_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({48885659, 205681680, 46120362, 175949223, 233437339, 127163336, 79843127, 90149574,
              158914825, 248133554, 264322432, 229032903, 7376627, 4643973, 120080647, 98269185,
              92379159, 160048836, 184522009, 254234203, 100343421, 195181845, 66412546, 126749676,
              247452694, 266777211, 12551837, 161345834, 255457916, 59214954, 110302060, 135080569}))
  stage_2_butterfly_26 (
    .x_in(stage_1_per_out[52]),
    .y_in(stage_1_per_out[53]),
    .x_out(stage_2_per_in[52]),
    .y_out(stage_2_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({48885659, 205681680, 46120362, 175949223, 233437339, 127163336, 79843127, 90149574,
              158914825, 248133554, 264322432, 229032903, 7376627, 4643973, 120080647, 98269185,
              92379159, 160048836, 184522009, 254234203, 100343421, 195181845, 66412546, 126749676,
              247452694, 266777211, 12551837, 161345834, 255457916, 59214954, 110302060, 135080569}))
  stage_2_butterfly_27 (
    .x_in(stage_1_per_out[54]),
    .y_in(stage_1_per_out[55]),
    .x_out(stage_2_per_in[54]),
    .y_out(stage_2_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({2017030, 166139329, 20118393, 112756762, 95713937, 224550271, 67209795, 248465751,
              216531417, 171841734, 10943590, 7280660, 267017218, 105443909, 154298223, 247116469,
              227628318, 138513718, 166586238, 75689102, 195298807, 266777383, 265028258, 151297332,
              228243008, 104290760, 67241659, 176972907, 116257755, 27298769, 122455193, 208475153}))
  stage_2_butterfly_28 (
    .x_in(stage_1_per_out[56]),
    .y_in(stage_1_per_out[57]),
    .x_out(stage_2_per_in[56]),
    .y_out(stage_2_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({2017030, 166139329, 20118393, 112756762, 95713937, 224550271, 67209795, 248465751,
              216531417, 171841734, 10943590, 7280660, 267017218, 105443909, 154298223, 247116469,
              227628318, 138513718, 166586238, 75689102, 195298807, 266777383, 265028258, 151297332,
              228243008, 104290760, 67241659, 176972907, 116257755, 27298769, 122455193, 208475153}))
  stage_2_butterfly_29 (
    .x_in(stage_1_per_out[58]),
    .y_in(stage_1_per_out[59]),
    .x_out(stage_2_per_in[58]),
    .y_out(stage_2_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({2017030, 166139329, 20118393, 112756762, 95713937, 224550271, 67209795, 248465751,
              216531417, 171841734, 10943590, 7280660, 267017218, 105443909, 154298223, 247116469,
              227628318, 138513718, 166586238, 75689102, 195298807, 266777383, 265028258, 151297332,
              228243008, 104290760, 67241659, 176972907, 116257755, 27298769, 122455193, 208475153}))
  stage_2_butterfly_30 (
    .x_in(stage_1_per_out[60]),
    .y_in(stage_1_per_out[61]),
    .x_out(stage_2_per_in[60]),
    .y_out(stage_2_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({2017030, 166139329, 20118393, 112756762, 95713937, 224550271, 67209795, 248465751,
              216531417, 171841734, 10943590, 7280660, 267017218, 105443909, 154298223, 247116469,
              227628318, 138513718, 166586238, 75689102, 195298807, 266777383, 265028258, 151297332,
              228243008, 104290760, 67241659, 176972907, 116257755, 27298769, 122455193, 208475153}))
  stage_2_butterfly_31 (
    .x_in(stage_1_per_out[62]),
    .y_in(stage_1_per_out[63]),
    .x_out(stage_2_per_in[62]),
    .y_out(stage_2_per_in[63]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({235273242, 135902522, 249576229, 122969043, 206341936, 81414740, 141956852, 209112367,
              72369588, 265348407, 1855205, 171206517, 226834391, 77127228, 43000087, 246787643,
              237125965, 244423105, 85740049, 90687088, 167645260, 145831337, 206116619, 191744986,
              121730405, 205856513, 174028560, 175598948, 4721397, 146344523, 62435894, 193174373}))
  stage_2_butterfly_32 (
    .x_in(stage_1_per_out[64]),
    .y_in(stage_1_per_out[65]),
    .x_out(stage_2_per_in[64]),
    .y_out(stage_2_per_in[65]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({235273242, 135902522, 249576229, 122969043, 206341936, 81414740, 141956852, 209112367,
              72369588, 265348407, 1855205, 171206517, 226834391, 77127228, 43000087, 246787643,
              237125965, 244423105, 85740049, 90687088, 167645260, 145831337, 206116619, 191744986,
              121730405, 205856513, 174028560, 175598948, 4721397, 146344523, 62435894, 193174373}))
  stage_2_butterfly_33 (
    .x_in(stage_1_per_out[66]),
    .y_in(stage_1_per_out[67]),
    .x_out(stage_2_per_in[66]),
    .y_out(stage_2_per_in[67]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({235273242, 135902522, 249576229, 122969043, 206341936, 81414740, 141956852, 209112367,
              72369588, 265348407, 1855205, 171206517, 226834391, 77127228, 43000087, 246787643,
              237125965, 244423105, 85740049, 90687088, 167645260, 145831337, 206116619, 191744986,
              121730405, 205856513, 174028560, 175598948, 4721397, 146344523, 62435894, 193174373}))
  stage_2_butterfly_34 (
    .x_in(stage_1_per_out[68]),
    .y_in(stage_1_per_out[69]),
    .x_out(stage_2_per_in[68]),
    .y_out(stage_2_per_in[69]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({235273242, 135902522, 249576229, 122969043, 206341936, 81414740, 141956852, 209112367,
              72369588, 265348407, 1855205, 171206517, 226834391, 77127228, 43000087, 246787643,
              237125965, 244423105, 85740049, 90687088, 167645260, 145831337, 206116619, 191744986,
              121730405, 205856513, 174028560, 175598948, 4721397, 146344523, 62435894, 193174373}))
  stage_2_butterfly_35 (
    .x_in(stage_1_per_out[70]),
    .y_in(stage_1_per_out[71]),
    .x_out(stage_2_per_in[70]),
    .y_out(stage_2_per_in[71]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({77536776, 189601976, 155363318, 94792077, 65889055, 164248031, 212237706, 261541195,
              205242220, 34052825, 86359417, 254842567, 169792793, 146205579, 256834872, 159538295,
              250727821, 243339369, 56723699, 224922683, 191250025, 136179523, 61322741, 57946842,
              100611174, 56545684, 148479452, 161217010, 141267184, 5739737, 223481427, 103896237}))
  stage_2_butterfly_36 (
    .x_in(stage_1_per_out[72]),
    .y_in(stage_1_per_out[73]),
    .x_out(stage_2_per_in[72]),
    .y_out(stage_2_per_in[73]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({77536776, 189601976, 155363318, 94792077, 65889055, 164248031, 212237706, 261541195,
              205242220, 34052825, 86359417, 254842567, 169792793, 146205579, 256834872, 159538295,
              250727821, 243339369, 56723699, 224922683, 191250025, 136179523, 61322741, 57946842,
              100611174, 56545684, 148479452, 161217010, 141267184, 5739737, 223481427, 103896237}))
  stage_2_butterfly_37 (
    .x_in(stage_1_per_out[74]),
    .y_in(stage_1_per_out[75]),
    .x_out(stage_2_per_in[74]),
    .y_out(stage_2_per_in[75]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({77536776, 189601976, 155363318, 94792077, 65889055, 164248031, 212237706, 261541195,
              205242220, 34052825, 86359417, 254842567, 169792793, 146205579, 256834872, 159538295,
              250727821, 243339369, 56723699, 224922683, 191250025, 136179523, 61322741, 57946842,
              100611174, 56545684, 148479452, 161217010, 141267184, 5739737, 223481427, 103896237}))
  stage_2_butterfly_38 (
    .x_in(stage_1_per_out[76]),
    .y_in(stage_1_per_out[77]),
    .x_out(stage_2_per_in[76]),
    .y_out(stage_2_per_in[77]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({77536776, 189601976, 155363318, 94792077, 65889055, 164248031, 212237706, 261541195,
              205242220, 34052825, 86359417, 254842567, 169792793, 146205579, 256834872, 159538295,
              250727821, 243339369, 56723699, 224922683, 191250025, 136179523, 61322741, 57946842,
              100611174, 56545684, 148479452, 161217010, 141267184, 5739737, 223481427, 103896237}))
  stage_2_butterfly_39 (
    .x_in(stage_1_per_out[78]),
    .y_in(stage_1_per_out[79]),
    .x_out(stage_2_per_in[78]),
    .y_out(stage_2_per_in[79]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({73481957, 116513948, 89028484, 187106042, 207877484, 58903295, 12286825, 77916555,
              181167176, 145351880, 160204962, 45355620, 129325164, 259302720, 51550886, 110378476,
              218380292, 140358303, 3260661, 19058782, 190540901, 222527593, 60600589, 202565947,
              50174239, 226759664, 46197346, 92902456, 78552959, 159148996, 76313029, 24036023}))
  stage_2_butterfly_40 (
    .x_in(stage_1_per_out[80]),
    .y_in(stage_1_per_out[81]),
    .x_out(stage_2_per_in[80]),
    .y_out(stage_2_per_in[81]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({73481957, 116513948, 89028484, 187106042, 207877484, 58903295, 12286825, 77916555,
              181167176, 145351880, 160204962, 45355620, 129325164, 259302720, 51550886, 110378476,
              218380292, 140358303, 3260661, 19058782, 190540901, 222527593, 60600589, 202565947,
              50174239, 226759664, 46197346, 92902456, 78552959, 159148996, 76313029, 24036023}))
  stage_2_butterfly_41 (
    .x_in(stage_1_per_out[82]),
    .y_in(stage_1_per_out[83]),
    .x_out(stage_2_per_in[82]),
    .y_out(stage_2_per_in[83]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({73481957, 116513948, 89028484, 187106042, 207877484, 58903295, 12286825, 77916555,
              181167176, 145351880, 160204962, 45355620, 129325164, 259302720, 51550886, 110378476,
              218380292, 140358303, 3260661, 19058782, 190540901, 222527593, 60600589, 202565947,
              50174239, 226759664, 46197346, 92902456, 78552959, 159148996, 76313029, 24036023}))
  stage_2_butterfly_42 (
    .x_in(stage_1_per_out[84]),
    .y_in(stage_1_per_out[85]),
    .x_out(stage_2_per_in[84]),
    .y_out(stage_2_per_in[85]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({73481957, 116513948, 89028484, 187106042, 207877484, 58903295, 12286825, 77916555,
              181167176, 145351880, 160204962, 45355620, 129325164, 259302720, 51550886, 110378476,
              218380292, 140358303, 3260661, 19058782, 190540901, 222527593, 60600589, 202565947,
              50174239, 226759664, 46197346, 92902456, 78552959, 159148996, 76313029, 24036023}))
  stage_2_butterfly_43 (
    .x_in(stage_1_per_out[86]),
    .y_in(stage_1_per_out[87]),
    .x_out(stage_2_per_in[86]),
    .y_out(stage_2_per_in[87]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({183700349, 188535281, 174391063, 266378632, 150049787, 189044804, 175710456, 104215821,
              159987098, 140210175, 72677507, 197425604, 92441360, 58726750, 236050384, 153319834,
              135921552, 161607031, 9793208, 52844710, 69205492, 187867192, 164728317, 243091016,
              8650362, 8259535, 79336225, 234786570, 123052007, 261458154, 129740611, 2204580}))
  stage_2_butterfly_44 (
    .x_in(stage_1_per_out[88]),
    .y_in(stage_1_per_out[89]),
    .x_out(stage_2_per_in[88]),
    .y_out(stage_2_per_in[89]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({183700349, 188535281, 174391063, 266378632, 150049787, 189044804, 175710456, 104215821,
              159987098, 140210175, 72677507, 197425604, 92441360, 58726750, 236050384, 153319834,
              135921552, 161607031, 9793208, 52844710, 69205492, 187867192, 164728317, 243091016,
              8650362, 8259535, 79336225, 234786570, 123052007, 261458154, 129740611, 2204580}))
  stage_2_butterfly_45 (
    .x_in(stage_1_per_out[90]),
    .y_in(stage_1_per_out[91]),
    .x_out(stage_2_per_in[90]),
    .y_out(stage_2_per_in[91]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({183700349, 188535281, 174391063, 266378632, 150049787, 189044804, 175710456, 104215821,
              159987098, 140210175, 72677507, 197425604, 92441360, 58726750, 236050384, 153319834,
              135921552, 161607031, 9793208, 52844710, 69205492, 187867192, 164728317, 243091016,
              8650362, 8259535, 79336225, 234786570, 123052007, 261458154, 129740611, 2204580}))
  stage_2_butterfly_46 (
    .x_in(stage_1_per_out[92]),
    .y_in(stage_1_per_out[93]),
    .x_out(stage_2_per_in[92]),
    .y_out(stage_2_per_in[93]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({183700349, 188535281, 174391063, 266378632, 150049787, 189044804, 175710456, 104215821,
              159987098, 140210175, 72677507, 197425604, 92441360, 58726750, 236050384, 153319834,
              135921552, 161607031, 9793208, 52844710, 69205492, 187867192, 164728317, 243091016,
              8650362, 8259535, 79336225, 234786570, 123052007, 261458154, 129740611, 2204580}))
  stage_2_butterfly_47 (
    .x_in(stage_1_per_out[94]),
    .y_in(stage_1_per_out[95]),
    .x_out(stage_2_per_in[94]),
    .y_out(stage_2_per_in[95]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({266562472, 232847226, 83977288, 144502563, 262112169, 107503597, 217359458, 184177651,
              172401093, 5161923, 22997488, 252018541, 584543, 183571221, 198336839, 66582189,
              142807968, 174290656, 87492030, 22383105, 46312994, 238775640, 248328138, 250611881,
              209698557, 227453822, 93513491, 169092523, 258059551, 139742686, 131659168, 113269084}))
  stage_2_butterfly_48 (
    .x_in(stage_1_per_out[96]),
    .y_in(stage_1_per_out[97]),
    .x_out(stage_2_per_in[96]),
    .y_out(stage_2_per_in[97]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({266562472, 232847226, 83977288, 144502563, 262112169, 107503597, 217359458, 184177651,
              172401093, 5161923, 22997488, 252018541, 584543, 183571221, 198336839, 66582189,
              142807968, 174290656, 87492030, 22383105, 46312994, 238775640, 248328138, 250611881,
              209698557, 227453822, 93513491, 169092523, 258059551, 139742686, 131659168, 113269084}))
  stage_2_butterfly_49 (
    .x_in(stage_1_per_out[98]),
    .y_in(stage_1_per_out[99]),
    .x_out(stage_2_per_in[98]),
    .y_out(stage_2_per_in[99]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({266562472, 232847226, 83977288, 144502563, 262112169, 107503597, 217359458, 184177651,
              172401093, 5161923, 22997488, 252018541, 584543, 183571221, 198336839, 66582189,
              142807968, 174290656, 87492030, 22383105, 46312994, 238775640, 248328138, 250611881,
              209698557, 227453822, 93513491, 169092523, 258059551, 139742686, 131659168, 113269084}))
  stage_2_butterfly_50 (
    .x_in(stage_1_per_out[100]),
    .y_in(stage_1_per_out[101]),
    .x_out(stage_2_per_in[100]),
    .y_out(stage_2_per_in[101]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({266562472, 232847226, 83977288, 144502563, 262112169, 107503597, 217359458, 184177651,
              172401093, 5161923, 22997488, 252018541, 584543, 183571221, 198336839, 66582189,
              142807968, 174290656, 87492030, 22383105, 46312994, 238775640, 248328138, 250611881,
              209698557, 227453822, 93513491, 169092523, 258059551, 139742686, 131659168, 113269084}))
  stage_2_butterfly_51 (
    .x_in(stage_1_per_out[102]),
    .y_in(stage_1_per_out[103]),
    .x_out(stage_2_per_in[102]),
    .y_out(stage_2_per_in[103]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({65498827, 181593250, 73685379, 133098101, 245041907, 133952844, 69412414, 149904904,
              265496406, 55947412, 134561032, 131471427, 228572460, 121970089, 186476418, 120318911,
              149925004, 236528116, 210373784, 53126225, 137060289, 255737752, 4457103, 157386503,
              23776027, 212162524, 203905228, 50376784, 203598031, 134804553, 193897399, 149423455}))
  stage_2_butterfly_52 (
    .x_in(stage_1_per_out[104]),
    .y_in(stage_1_per_out[105]),
    .x_out(stage_2_per_in[104]),
    .y_out(stage_2_per_in[105]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({65498827, 181593250, 73685379, 133098101, 245041907, 133952844, 69412414, 149904904,
              265496406, 55947412, 134561032, 131471427, 228572460, 121970089, 186476418, 120318911,
              149925004, 236528116, 210373784, 53126225, 137060289, 255737752, 4457103, 157386503,
              23776027, 212162524, 203905228, 50376784, 203598031, 134804553, 193897399, 149423455}))
  stage_2_butterfly_53 (
    .x_in(stage_1_per_out[106]),
    .y_in(stage_1_per_out[107]),
    .x_out(stage_2_per_in[106]),
    .y_out(stage_2_per_in[107]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({65498827, 181593250, 73685379, 133098101, 245041907, 133952844, 69412414, 149904904,
              265496406, 55947412, 134561032, 131471427, 228572460, 121970089, 186476418, 120318911,
              149925004, 236528116, 210373784, 53126225, 137060289, 255737752, 4457103, 157386503,
              23776027, 212162524, 203905228, 50376784, 203598031, 134804553, 193897399, 149423455}))
  stage_2_butterfly_54 (
    .x_in(stage_1_per_out[108]),
    .y_in(stage_1_per_out[109]),
    .x_out(stage_2_per_in[108]),
    .y_out(stage_2_per_in[109]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({65498827, 181593250, 73685379, 133098101, 245041907, 133952844, 69412414, 149904904,
              265496406, 55947412, 134561032, 131471427, 228572460, 121970089, 186476418, 120318911,
              149925004, 236528116, 210373784, 53126225, 137060289, 255737752, 4457103, 157386503,
              23776027, 212162524, 203905228, 50376784, 203598031, 134804553, 193897399, 149423455}))
  stage_2_butterfly_55 (
    .x_in(stage_1_per_out[110]),
    .y_in(stage_1_per_out[111]),
    .x_out(stage_2_per_in[110]),
    .y_out(stage_2_per_in[111]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({98410858, 16697663, 163823140, 56081948, 121712648, 53432143, 265883664, 94856770,
              126807666, 23586243, 123313741, 232038388, 217846048, 106743034, 121145061, 2487567,
              6001670, 55581691, 170230234, 180764097, 103503994, 37498403, 99996719, 5445105,
              62094530, 219133933, 55222727, 183669067, 263649093, 101579460, 7301415, 168342750}))
  stage_2_butterfly_56 (
    .x_in(stage_1_per_out[112]),
    .y_in(stage_1_per_out[113]),
    .x_out(stage_2_per_in[112]),
    .y_out(stage_2_per_in[113]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({98410858, 16697663, 163823140, 56081948, 121712648, 53432143, 265883664, 94856770,
              126807666, 23586243, 123313741, 232038388, 217846048, 106743034, 121145061, 2487567,
              6001670, 55581691, 170230234, 180764097, 103503994, 37498403, 99996719, 5445105,
              62094530, 219133933, 55222727, 183669067, 263649093, 101579460, 7301415, 168342750}))
  stage_2_butterfly_57 (
    .x_in(stage_1_per_out[114]),
    .y_in(stage_1_per_out[115]),
    .x_out(stage_2_per_in[114]),
    .y_out(stage_2_per_in[115]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({98410858, 16697663, 163823140, 56081948, 121712648, 53432143, 265883664, 94856770,
              126807666, 23586243, 123313741, 232038388, 217846048, 106743034, 121145061, 2487567,
              6001670, 55581691, 170230234, 180764097, 103503994, 37498403, 99996719, 5445105,
              62094530, 219133933, 55222727, 183669067, 263649093, 101579460, 7301415, 168342750}))
  stage_2_butterfly_58 (
    .x_in(stage_1_per_out[116]),
    .y_in(stage_1_per_out[117]),
    .x_out(stage_2_per_in[116]),
    .y_out(stage_2_per_in[117]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({98410858, 16697663, 163823140, 56081948, 121712648, 53432143, 265883664, 94856770,
              126807666, 23586243, 123313741, 232038388, 217846048, 106743034, 121145061, 2487567,
              6001670, 55581691, 170230234, 180764097, 103503994, 37498403, 99996719, 5445105,
              62094530, 219133933, 55222727, 183669067, 263649093, 101579460, 7301415, 168342750}))
  stage_2_butterfly_59 (
    .x_in(stage_1_per_out[118]),
    .y_in(stage_1_per_out[119]),
    .x_out(stage_2_per_in[118]),
    .y_out(stage_2_per_in[119]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({217210388, 17682401, 60051251, 107138937, 209744644, 86350556, 112825183, 24347842,
              62765404, 19637177, 81197166, 244216061, 223473865, 29901564, 160429892, 30998914,
              102243739, 21628090, 226981541, 95654178, 198352904, 189248215, 103189081, 231749609,
              58589536, 74931497, 255778637, 178382895, 80381167, 203850982, 18433789, 98445813}))
  stage_2_butterfly_60 (
    .x_in(stage_1_per_out[120]),
    .y_in(stage_1_per_out[121]),
    .x_out(stage_2_per_in[120]),
    .y_out(stage_2_per_in[121]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({217210388, 17682401, 60051251, 107138937, 209744644, 86350556, 112825183, 24347842,
              62765404, 19637177, 81197166, 244216061, 223473865, 29901564, 160429892, 30998914,
              102243739, 21628090, 226981541, 95654178, 198352904, 189248215, 103189081, 231749609,
              58589536, 74931497, 255778637, 178382895, 80381167, 203850982, 18433789, 98445813}))
  stage_2_butterfly_61 (
    .x_in(stage_1_per_out[122]),
    .y_in(stage_1_per_out[123]),
    .x_out(stage_2_per_in[122]),
    .y_out(stage_2_per_in[123]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({217210388, 17682401, 60051251, 107138937, 209744644, 86350556, 112825183, 24347842,
              62765404, 19637177, 81197166, 244216061, 223473865, 29901564, 160429892, 30998914,
              102243739, 21628090, 226981541, 95654178, 198352904, 189248215, 103189081, 231749609,
              58589536, 74931497, 255778637, 178382895, 80381167, 203850982, 18433789, 98445813}))
  stage_2_butterfly_62 (
    .x_in(stage_1_per_out[124]),
    .y_in(stage_1_per_out[125]),
    .x_out(stage_2_per_in[124]),
    .y_out(stage_2_per_in[125]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({217210388, 17682401, 60051251, 107138937, 209744644, 86350556, 112825183, 24347842,
              62765404, 19637177, 81197166, 244216061, 223473865, 29901564, 160429892, 30998914,
              102243739, 21628090, 226981541, 95654178, 198352904, 189248215, 103189081, 231749609,
              58589536, 74931497, 255778637, 178382895, 80381167, 203850982, 18433789, 98445813}))
  stage_2_butterfly_63 (
    .x_in(stage_1_per_out[126]),
    .y_in(stage_1_per_out[127]),
    .x_out(stage_2_per_in[126]),
    .y_out(stage_2_per_in[127]),
    .clk(clk),
    .rst(rst)
  );



  // TODO(Yang): stage 2 -> stage 3 permutation
  // FIXME: ignore butterfly units for now.
  stage_2_permutation #(
    .DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    .INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_2_3_per (
    .inData_0(stage_2_per_in[0]),
    .inData_1(stage_2_per_in[1]),
    .inData_2(stage_2_per_in[2]),
    .inData_3(stage_2_per_in[3]),
    .inData_4(stage_2_per_in[4]),
    .inData_5(stage_2_per_in[5]),
    .inData_6(stage_2_per_in[6]),
    .inData_7(stage_2_per_in[7]),
    .inData_8(stage_2_per_in[8]),
    .inData_9(stage_2_per_in[9]),
    .inData_10(stage_2_per_in[10]),
    .inData_11(stage_2_per_in[11]),
    .inData_12(stage_2_per_in[12]),
    .inData_13(stage_2_per_in[13]),
    .inData_14(stage_2_per_in[14]),
    .inData_15(stage_2_per_in[15]),
    .inData_16(stage_2_per_in[16]),
    .inData_17(stage_2_per_in[17]),
    .inData_18(stage_2_per_in[18]),
    .inData_19(stage_2_per_in[19]),
    .inData_20(stage_2_per_in[20]),
    .inData_21(stage_2_per_in[21]),
    .inData_22(stage_2_per_in[22]),
    .inData_23(stage_2_per_in[23]),
    .inData_24(stage_2_per_in[24]),
    .inData_25(stage_2_per_in[25]),
    .inData_26(stage_2_per_in[26]),
    .inData_27(stage_2_per_in[27]),
    .inData_28(stage_2_per_in[28]),
    .inData_29(stage_2_per_in[29]),
    .inData_30(stage_2_per_in[30]),
    .inData_31(stage_2_per_in[31]),
    .inData_32(stage_2_per_in[32]),
    .inData_33(stage_2_per_in[33]),
    .inData_34(stage_2_per_in[34]),
    .inData_35(stage_2_per_in[35]),
    .inData_36(stage_2_per_in[36]),
    .inData_37(stage_2_per_in[37]),
    .inData_38(stage_2_per_in[38]),
    .inData_39(stage_2_per_in[39]),
    .inData_40(stage_2_per_in[40]),
    .inData_41(stage_2_per_in[41]),
    .inData_42(stage_2_per_in[42]),
    .inData_43(stage_2_per_in[43]),
    .inData_44(stage_2_per_in[44]),
    .inData_45(stage_2_per_in[45]),
    .inData_46(stage_2_per_in[46]),
    .inData_47(stage_2_per_in[47]),
    .inData_48(stage_2_per_in[48]),
    .inData_49(stage_2_per_in[49]),
    .inData_50(stage_2_per_in[50]),
    .inData_51(stage_2_per_in[51]),
    .inData_52(stage_2_per_in[52]),
    .inData_53(stage_2_per_in[53]),
    .inData_54(stage_2_per_in[54]),
    .inData_55(stage_2_per_in[55]),
    .inData_56(stage_2_per_in[56]),
    .inData_57(stage_2_per_in[57]),
    .inData_58(stage_2_per_in[58]),
    .inData_59(stage_2_per_in[59]),
    .inData_60(stage_2_per_in[60]),
    .inData_61(stage_2_per_in[61]),
    .inData_62(stage_2_per_in[62]),
    .inData_63(stage_2_per_in[63]),
    .inData_64(stage_2_per_in[64]),
    .inData_65(stage_2_per_in[65]),
    .inData_66(stage_2_per_in[66]),
    .inData_67(stage_2_per_in[67]),
    .inData_68(stage_2_per_in[68]),
    .inData_69(stage_2_per_in[69]),
    .inData_70(stage_2_per_in[70]),
    .inData_71(stage_2_per_in[71]),
    .inData_72(stage_2_per_in[72]),
    .inData_73(stage_2_per_in[73]),
    .inData_74(stage_2_per_in[74]),
    .inData_75(stage_2_per_in[75]),
    .inData_76(stage_2_per_in[76]),
    .inData_77(stage_2_per_in[77]),
    .inData_78(stage_2_per_in[78]),
    .inData_79(stage_2_per_in[79]),
    .inData_80(stage_2_per_in[80]),
    .inData_81(stage_2_per_in[81]),
    .inData_82(stage_2_per_in[82]),
    .inData_83(stage_2_per_in[83]),
    .inData_84(stage_2_per_in[84]),
    .inData_85(stage_2_per_in[85]),
    .inData_86(stage_2_per_in[86]),
    .inData_87(stage_2_per_in[87]),
    .inData_88(stage_2_per_in[88]),
    .inData_89(stage_2_per_in[89]),
    .inData_90(stage_2_per_in[90]),
    .inData_91(stage_2_per_in[91]),
    .inData_92(stage_2_per_in[92]),
    .inData_93(stage_2_per_in[93]),
    .inData_94(stage_2_per_in[94]),
    .inData_95(stage_2_per_in[95]),
    .inData_96(stage_2_per_in[96]),
    .inData_97(stage_2_per_in[97]),
    .inData_98(stage_2_per_in[98]),
    .inData_99(stage_2_per_in[99]),
    .inData_100(stage_2_per_in[100]),
    .inData_101(stage_2_per_in[101]),
    .inData_102(stage_2_per_in[102]),
    .inData_103(stage_2_per_in[103]),
    .inData_104(stage_2_per_in[104]),
    .inData_105(stage_2_per_in[105]),
    .inData_106(stage_2_per_in[106]),
    .inData_107(stage_2_per_in[107]),
    .inData_108(stage_2_per_in[108]),
    .inData_109(stage_2_per_in[109]),
    .inData_110(stage_2_per_in[110]),
    .inData_111(stage_2_per_in[111]),
    .inData_112(stage_2_per_in[112]),
    .inData_113(stage_2_per_in[113]),
    .inData_114(stage_2_per_in[114]),
    .inData_115(stage_2_per_in[115]),
    .inData_116(stage_2_per_in[116]),
    .inData_117(stage_2_per_in[117]),
    .inData_118(stage_2_per_in[118]),
    .inData_119(stage_2_per_in[119]),
    .inData_120(stage_2_per_in[120]),
    .inData_121(stage_2_per_in[121]),
    .inData_122(stage_2_per_in[122]),
    .inData_123(stage_2_per_in[123]),
    .inData_124(stage_2_per_in[124]),
    .inData_125(stage_2_per_in[125]),
    .inData_126(stage_2_per_in[126]),
    .inData_127(stage_2_per_in[127]),
    .outData_0(stage_2_per_out[0]),
    .outData_1(stage_2_per_out[1]),
    .outData_2(stage_2_per_out[2]),
    .outData_3(stage_2_per_out[3]),
    .outData_4(stage_2_per_out[4]),
    .outData_5(stage_2_per_out[5]),
    .outData_6(stage_2_per_out[6]),
    .outData_7(stage_2_per_out[7]),
    .outData_8(stage_2_per_out[8]),
    .outData_9(stage_2_per_out[9]),
    .outData_10(stage_2_per_out[10]),
    .outData_11(stage_2_per_out[11]),
    .outData_12(stage_2_per_out[12]),
    .outData_13(stage_2_per_out[13]),
    .outData_14(stage_2_per_out[14]),
    .outData_15(stage_2_per_out[15]),
    .outData_16(stage_2_per_out[16]),
    .outData_17(stage_2_per_out[17]),
    .outData_18(stage_2_per_out[18]),
    .outData_19(stage_2_per_out[19]),
    .outData_20(stage_2_per_out[20]),
    .outData_21(stage_2_per_out[21]),
    .outData_22(stage_2_per_out[22]),
    .outData_23(stage_2_per_out[23]),
    .outData_24(stage_2_per_out[24]),
    .outData_25(stage_2_per_out[25]),
    .outData_26(stage_2_per_out[26]),
    .outData_27(stage_2_per_out[27]),
    .outData_28(stage_2_per_out[28]),
    .outData_29(stage_2_per_out[29]),
    .outData_30(stage_2_per_out[30]),
    .outData_31(stage_2_per_out[31]),
    .outData_32(stage_2_per_out[32]),
    .outData_33(stage_2_per_out[33]),
    .outData_34(stage_2_per_out[34]),
    .outData_35(stage_2_per_out[35]),
    .outData_36(stage_2_per_out[36]),
    .outData_37(stage_2_per_out[37]),
    .outData_38(stage_2_per_out[38]),
    .outData_39(stage_2_per_out[39]),
    .outData_40(stage_2_per_out[40]),
    .outData_41(stage_2_per_out[41]),
    .outData_42(stage_2_per_out[42]),
    .outData_43(stage_2_per_out[43]),
    .outData_44(stage_2_per_out[44]),
    .outData_45(stage_2_per_out[45]),
    .outData_46(stage_2_per_out[46]),
    .outData_47(stage_2_per_out[47]),
    .outData_48(stage_2_per_out[48]),
    .outData_49(stage_2_per_out[49]),
    .outData_50(stage_2_per_out[50]),
    .outData_51(stage_2_per_out[51]),
    .outData_52(stage_2_per_out[52]),
    .outData_53(stage_2_per_out[53]),
    .outData_54(stage_2_per_out[54]),
    .outData_55(stage_2_per_out[55]),
    .outData_56(stage_2_per_out[56]),
    .outData_57(stage_2_per_out[57]),
    .outData_58(stage_2_per_out[58]),
    .outData_59(stage_2_per_out[59]),
    .outData_60(stage_2_per_out[60]),
    .outData_61(stage_2_per_out[61]),
    .outData_62(stage_2_per_out[62]),
    .outData_63(stage_2_per_out[63]),
    .outData_64(stage_2_per_out[64]),
    .outData_65(stage_2_per_out[65]),
    .outData_66(stage_2_per_out[66]),
    .outData_67(stage_2_per_out[67]),
    .outData_68(stage_2_per_out[68]),
    .outData_69(stage_2_per_out[69]),
    .outData_70(stage_2_per_out[70]),
    .outData_71(stage_2_per_out[71]),
    .outData_72(stage_2_per_out[72]),
    .outData_73(stage_2_per_out[73]),
    .outData_74(stage_2_per_out[74]),
    .outData_75(stage_2_per_out[75]),
    .outData_76(stage_2_per_out[76]),
    .outData_77(stage_2_per_out[77]),
    .outData_78(stage_2_per_out[78]),
    .outData_79(stage_2_per_out[79]),
    .outData_80(stage_2_per_out[80]),
    .outData_81(stage_2_per_out[81]),
    .outData_82(stage_2_per_out[82]),
    .outData_83(stage_2_per_out[83]),
    .outData_84(stage_2_per_out[84]),
    .outData_85(stage_2_per_out[85]),
    .outData_86(stage_2_per_out[86]),
    .outData_87(stage_2_per_out[87]),
    .outData_88(stage_2_per_out[88]),
    .outData_89(stage_2_per_out[89]),
    .outData_90(stage_2_per_out[90]),
    .outData_91(stage_2_per_out[91]),
    .outData_92(stage_2_per_out[92]),
    .outData_93(stage_2_per_out[93]),
    .outData_94(stage_2_per_out[94]),
    .outData_95(stage_2_per_out[95]),
    .outData_96(stage_2_per_out[96]),
    .outData_97(stage_2_per_out[97]),
    .outData_98(stage_2_per_out[98]),
    .outData_99(stage_2_per_out[99]),
    .outData_100(stage_2_per_out[100]),
    .outData_101(stage_2_per_out[101]),
    .outData_102(stage_2_per_out[102]),
    .outData_103(stage_2_per_out[103]),
    .outData_104(stage_2_per_out[104]),
    .outData_105(stage_2_per_out[105]),
    .outData_106(stage_2_per_out[106]),
    .outData_107(stage_2_per_out[107]),
    .outData_108(stage_2_per_out[108]),
    .outData_109(stage_2_per_out[109]),
    .outData_110(stage_2_per_out[110]),
    .outData_111(stage_2_per_out[111]),
    .outData_112(stage_2_per_out[112]),
    .outData_113(stage_2_per_out[113]),
    .outData_114(stage_2_per_out[114]),
    .outData_115(stage_2_per_out[115]),
    .outData_116(stage_2_per_out[116]),
    .outData_117(stage_2_per_out[117]),
    .outData_118(stage_2_per_out[118]),
    .outData_119(stage_2_per_out[119]),
    .outData_120(stage_2_per_out[120]),
    .outData_121(stage_2_per_out[121]),
    .outData_122(stage_2_per_out[122]),
    .outData_123(stage_2_per_out[123]),
    .outData_124(stage_2_per_out[124]),
    .outData_125(stage_2_per_out[125]),
    .outData_126(stage_2_per_out[126]),
    .outData_127(stage_2_per_out[127]),
    .in_start(in_start[2]),
    .out_start(out_start[2]),
    .clk(clk),
    .rst(rst)
  );

  // TODO(Tian): stage 3 32 butterfly units
  butterfly #(
    .start(START_CYCLE[3]),
    .factors({135618975, 141849606, 98889920, 134877507, 64884498, 186863562, 224068691, 100123291,
              209658551, 99392088, 258527796, 85252512, 65324949, 95282463, 227819465, 20857483,
              198785423, 1562592, 219083512, 194276347, 251898247, 44144526, 255286072, 170930026,
              224794776, 176665584, 202776751, 246630386, 165872957, 172508742, 73698550, 208297913}))
  stage_3_butterfly_0 (
    .x_in(stage_2_per_out[0]),
    .y_in(stage_2_per_out[1]),
    .x_out(stage_3_per_in[0]),
    .y_out(stage_3_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({135618975, 141849606, 98889920, 134877507, 64884498, 186863562, 224068691, 100123291,
              209658551, 99392088, 258527796, 85252512, 65324949, 95282463, 227819465, 20857483,
              198785423, 1562592, 219083512, 194276347, 251898247, 44144526, 255286072, 170930026,
              224794776, 176665584, 202776751, 246630386, 165872957, 172508742, 73698550, 208297913}))
  stage_3_butterfly_1 (
    .x_in(stage_2_per_out[2]),
    .y_in(stage_2_per_out[3]),
    .x_out(stage_3_per_in[2]),
    .y_out(stage_3_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({135618975, 141849606, 98889920, 134877507, 64884498, 186863562, 224068691, 100123291,
              209658551, 99392088, 258527796, 85252512, 65324949, 95282463, 227819465, 20857483,
              198785423, 1562592, 219083512, 194276347, 251898247, 44144526, 255286072, 170930026,
              224794776, 176665584, 202776751, 246630386, 165872957, 172508742, 73698550, 208297913}))
  stage_3_butterfly_2 (
    .x_in(stage_2_per_out[4]),
    .y_in(stage_2_per_out[5]),
    .x_out(stage_3_per_in[4]),
    .y_out(stage_3_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({135618975, 141849606, 98889920, 134877507, 64884498, 186863562, 224068691, 100123291,
              209658551, 99392088, 258527796, 85252512, 65324949, 95282463, 227819465, 20857483,
              198785423, 1562592, 219083512, 194276347, 251898247, 44144526, 255286072, 170930026,
              224794776, 176665584, 202776751, 246630386, 165872957, 172508742, 73698550, 208297913}))
  stage_3_butterfly_3 (
    .x_in(stage_2_per_out[6]),
    .y_in(stage_2_per_out[7]),
    .x_out(stage_3_per_in[6]),
    .y_out(stage_3_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({135618975, 141849606, 98889920, 134877507, 64884498, 186863562, 224068691, 100123291,
              209658551, 99392088, 258527796, 85252512, 65324949, 95282463, 227819465, 20857483,
              198785423, 1562592, 219083512, 194276347, 251898247, 44144526, 255286072, 170930026,
              224794776, 176665584, 202776751, 246630386, 165872957, 172508742, 73698550, 208297913}))
  stage_3_butterfly_4 (
    .x_in(stage_2_per_out[8]),
    .y_in(stage_2_per_out[9]),
    .x_out(stage_3_per_in[8]),
    .y_out(stage_3_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({135618975, 141849606, 98889920, 134877507, 64884498, 186863562, 224068691, 100123291,
              209658551, 99392088, 258527796, 85252512, 65324949, 95282463, 227819465, 20857483,
              198785423, 1562592, 219083512, 194276347, 251898247, 44144526, 255286072, 170930026,
              224794776, 176665584, 202776751, 246630386, 165872957, 172508742, 73698550, 208297913}))
  stage_3_butterfly_5 (
    .x_in(stage_2_per_out[10]),
    .y_in(stage_2_per_out[11]),
    .x_out(stage_3_per_in[10]),
    .y_out(stage_3_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({135618975, 141849606, 98889920, 134877507, 64884498, 186863562, 224068691, 100123291,
              209658551, 99392088, 258527796, 85252512, 65324949, 95282463, 227819465, 20857483,
              198785423, 1562592, 219083512, 194276347, 251898247, 44144526, 255286072, 170930026,
              224794776, 176665584, 202776751, 246630386, 165872957, 172508742, 73698550, 208297913}))
  stage_3_butterfly_6 (
    .x_in(stage_2_per_out[12]),
    .y_in(stage_2_per_out[13]),
    .x_out(stage_3_per_in[12]),
    .y_out(stage_3_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({135618975, 141849606, 98889920, 134877507, 64884498, 186863562, 224068691, 100123291,
              209658551, 99392088, 258527796, 85252512, 65324949, 95282463, 227819465, 20857483,
              198785423, 1562592, 219083512, 194276347, 251898247, 44144526, 255286072, 170930026,
              224794776, 176665584, 202776751, 246630386, 165872957, 172508742, 73698550, 208297913}))
  stage_3_butterfly_7 (
    .x_in(stage_2_per_out[14]),
    .y_in(stage_2_per_out[15]),
    .x_out(stage_3_per_in[14]),
    .y_out(stage_3_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({42355602, 45686070, 78649100, 17861009, 160254284, 57574719, 117221766, 182702557,
              136878682, 5829490, 61345534, 148801771, 69773246, 56155754, 137065607, 40158424,
              54534442, 249146534, 61720173, 64764693, 258559590, 134269022, 184644727, 142306631,
              220994759, 8950678, 225784463, 61664240, 23892097, 234350511, 49504466, 66505970}))
  stage_3_butterfly_8 (
    .x_in(stage_2_per_out[16]),
    .y_in(stage_2_per_out[17]),
    .x_out(stage_3_per_in[16]),
    .y_out(stage_3_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({42355602, 45686070, 78649100, 17861009, 160254284, 57574719, 117221766, 182702557,
              136878682, 5829490, 61345534, 148801771, 69773246, 56155754, 137065607, 40158424,
              54534442, 249146534, 61720173, 64764693, 258559590, 134269022, 184644727, 142306631,
              220994759, 8950678, 225784463, 61664240, 23892097, 234350511, 49504466, 66505970}))
  stage_3_butterfly_9 (
    .x_in(stage_2_per_out[18]),
    .y_in(stage_2_per_out[19]),
    .x_out(stage_3_per_in[18]),
    .y_out(stage_3_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({42355602, 45686070, 78649100, 17861009, 160254284, 57574719, 117221766, 182702557,
              136878682, 5829490, 61345534, 148801771, 69773246, 56155754, 137065607, 40158424,
              54534442, 249146534, 61720173, 64764693, 258559590, 134269022, 184644727, 142306631,
              220994759, 8950678, 225784463, 61664240, 23892097, 234350511, 49504466, 66505970}))
  stage_3_butterfly_10 (
    .x_in(stage_2_per_out[20]),
    .y_in(stage_2_per_out[21]),
    .x_out(stage_3_per_in[20]),
    .y_out(stage_3_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({42355602, 45686070, 78649100, 17861009, 160254284, 57574719, 117221766, 182702557,
              136878682, 5829490, 61345534, 148801771, 69773246, 56155754, 137065607, 40158424,
              54534442, 249146534, 61720173, 64764693, 258559590, 134269022, 184644727, 142306631,
              220994759, 8950678, 225784463, 61664240, 23892097, 234350511, 49504466, 66505970}))
  stage_3_butterfly_11 (
    .x_in(stage_2_per_out[22]),
    .y_in(stage_2_per_out[23]),
    .x_out(stage_3_per_in[22]),
    .y_out(stage_3_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({42355602, 45686070, 78649100, 17861009, 160254284, 57574719, 117221766, 182702557,
              136878682, 5829490, 61345534, 148801771, 69773246, 56155754, 137065607, 40158424,
              54534442, 249146534, 61720173, 64764693, 258559590, 134269022, 184644727, 142306631,
              220994759, 8950678, 225784463, 61664240, 23892097, 234350511, 49504466, 66505970}))
  stage_3_butterfly_12 (
    .x_in(stage_2_per_out[24]),
    .y_in(stage_2_per_out[25]),
    .x_out(stage_3_per_in[24]),
    .y_out(stage_3_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({42355602, 45686070, 78649100, 17861009, 160254284, 57574719, 117221766, 182702557,
              136878682, 5829490, 61345534, 148801771, 69773246, 56155754, 137065607, 40158424,
              54534442, 249146534, 61720173, 64764693, 258559590, 134269022, 184644727, 142306631,
              220994759, 8950678, 225784463, 61664240, 23892097, 234350511, 49504466, 66505970}))
  stage_3_butterfly_13 (
    .x_in(stage_2_per_out[26]),
    .y_in(stage_2_per_out[27]),
    .x_out(stage_3_per_in[26]),
    .y_out(stage_3_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({42355602, 45686070, 78649100, 17861009, 160254284, 57574719, 117221766, 182702557,
              136878682, 5829490, 61345534, 148801771, 69773246, 56155754, 137065607, 40158424,
              54534442, 249146534, 61720173, 64764693, 258559590, 134269022, 184644727, 142306631,
              220994759, 8950678, 225784463, 61664240, 23892097, 234350511, 49504466, 66505970}))
  stage_3_butterfly_14 (
    .x_in(stage_2_per_out[28]),
    .y_in(stage_2_per_out[29]),
    .x_out(stage_3_per_in[28]),
    .y_out(stage_3_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({42355602, 45686070, 78649100, 17861009, 160254284, 57574719, 117221766, 182702557,
              136878682, 5829490, 61345534, 148801771, 69773246, 56155754, 137065607, 40158424,
              54534442, 249146534, 61720173, 64764693, 258559590, 134269022, 184644727, 142306631,
              220994759, 8950678, 225784463, 61664240, 23892097, 234350511, 49504466, 66505970}))
  stage_3_butterfly_15 (
    .x_in(stage_2_per_out[30]),
    .y_in(stage_2_per_out[31]),
    .x_out(stage_3_per_in[30]),
    .y_out(stage_3_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({98861208, 12196542, 232615475, 201144768, 253800975, 181295312, 205961920, 23606744,
              79852752, 32087335, 141424302, 172809179, 123440080, 94612904, 181468172, 16985430,
              233514072, 185685569, 172935357, 44547301, 93740850, 143102859, 109902969, 164638888,
              87202272, 57455860, 150862394, 161171966, 1613379, 6010959, 225291788, 215146927}))
  stage_3_butterfly_16 (
    .x_in(stage_2_per_out[32]),
    .y_in(stage_2_per_out[33]),
    .x_out(stage_3_per_in[32]),
    .y_out(stage_3_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({98861208, 12196542, 232615475, 201144768, 253800975, 181295312, 205961920, 23606744,
              79852752, 32087335, 141424302, 172809179, 123440080, 94612904, 181468172, 16985430,
              233514072, 185685569, 172935357, 44547301, 93740850, 143102859, 109902969, 164638888,
              87202272, 57455860, 150862394, 161171966, 1613379, 6010959, 225291788, 215146927}))
  stage_3_butterfly_17 (
    .x_in(stage_2_per_out[34]),
    .y_in(stage_2_per_out[35]),
    .x_out(stage_3_per_in[34]),
    .y_out(stage_3_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({98861208, 12196542, 232615475, 201144768, 253800975, 181295312, 205961920, 23606744,
              79852752, 32087335, 141424302, 172809179, 123440080, 94612904, 181468172, 16985430,
              233514072, 185685569, 172935357, 44547301, 93740850, 143102859, 109902969, 164638888,
              87202272, 57455860, 150862394, 161171966, 1613379, 6010959, 225291788, 215146927}))
  stage_3_butterfly_18 (
    .x_in(stage_2_per_out[36]),
    .y_in(stage_2_per_out[37]),
    .x_out(stage_3_per_in[36]),
    .y_out(stage_3_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({98861208, 12196542, 232615475, 201144768, 253800975, 181295312, 205961920, 23606744,
              79852752, 32087335, 141424302, 172809179, 123440080, 94612904, 181468172, 16985430,
              233514072, 185685569, 172935357, 44547301, 93740850, 143102859, 109902969, 164638888,
              87202272, 57455860, 150862394, 161171966, 1613379, 6010959, 225291788, 215146927}))
  stage_3_butterfly_19 (
    .x_in(stage_2_per_out[38]),
    .y_in(stage_2_per_out[39]),
    .x_out(stage_3_per_in[38]),
    .y_out(stage_3_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({98861208, 12196542, 232615475, 201144768, 253800975, 181295312, 205961920, 23606744,
              79852752, 32087335, 141424302, 172809179, 123440080, 94612904, 181468172, 16985430,
              233514072, 185685569, 172935357, 44547301, 93740850, 143102859, 109902969, 164638888,
              87202272, 57455860, 150862394, 161171966, 1613379, 6010959, 225291788, 215146927}))
  stage_3_butterfly_20 (
    .x_in(stage_2_per_out[40]),
    .y_in(stage_2_per_out[41]),
    .x_out(stage_3_per_in[40]),
    .y_out(stage_3_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({98861208, 12196542, 232615475, 201144768, 253800975, 181295312, 205961920, 23606744,
              79852752, 32087335, 141424302, 172809179, 123440080, 94612904, 181468172, 16985430,
              233514072, 185685569, 172935357, 44547301, 93740850, 143102859, 109902969, 164638888,
              87202272, 57455860, 150862394, 161171966, 1613379, 6010959, 225291788, 215146927}))
  stage_3_butterfly_21 (
    .x_in(stage_2_per_out[42]),
    .y_in(stage_2_per_out[43]),
    .x_out(stage_3_per_in[42]),
    .y_out(stage_3_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({98861208, 12196542, 232615475, 201144768, 253800975, 181295312, 205961920, 23606744,
              79852752, 32087335, 141424302, 172809179, 123440080, 94612904, 181468172, 16985430,
              233514072, 185685569, 172935357, 44547301, 93740850, 143102859, 109902969, 164638888,
              87202272, 57455860, 150862394, 161171966, 1613379, 6010959, 225291788, 215146927}))
  stage_3_butterfly_22 (
    .x_in(stage_2_per_out[44]),
    .y_in(stage_2_per_out[45]),
    .x_out(stage_3_per_in[44]),
    .y_out(stage_3_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({98861208, 12196542, 232615475, 201144768, 253800975, 181295312, 205961920, 23606744,
              79852752, 32087335, 141424302, 172809179, 123440080, 94612904, 181468172, 16985430,
              233514072, 185685569, 172935357, 44547301, 93740850, 143102859, 109902969, 164638888,
              87202272, 57455860, 150862394, 161171966, 1613379, 6010959, 225291788, 215146927}))
  stage_3_butterfly_23 (
    .x_in(stage_2_per_out[46]),
    .y_in(stage_2_per_out[47]),
    .x_out(stage_3_per_in[46]),
    .y_out(stage_3_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({77981460, 199633043, 142181410, 160841949, 8411857, 100229847, 75073484, 13458851,
              192832423, 56246211, 62117518, 148390399, 209085090, 10003248, 241313184, 25944135,
              212802310, 50222736, 18298478, 209886001, 145034471, 186841927, 160807241, 258257144,
              193915204, 92650808, 171362072, 30930936, 158727274, 226213489, 244216783, 158168844}))
  stage_3_butterfly_24 (
    .x_in(stage_2_per_out[48]),
    .y_in(stage_2_per_out[49]),
    .x_out(stage_3_per_in[48]),
    .y_out(stage_3_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({77981460, 199633043, 142181410, 160841949, 8411857, 100229847, 75073484, 13458851,
              192832423, 56246211, 62117518, 148390399, 209085090, 10003248, 241313184, 25944135,
              212802310, 50222736, 18298478, 209886001, 145034471, 186841927, 160807241, 258257144,
              193915204, 92650808, 171362072, 30930936, 158727274, 226213489, 244216783, 158168844}))
  stage_3_butterfly_25 (
    .x_in(stage_2_per_out[50]),
    .y_in(stage_2_per_out[51]),
    .x_out(stage_3_per_in[50]),
    .y_out(stage_3_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({77981460, 199633043, 142181410, 160841949, 8411857, 100229847, 75073484, 13458851,
              192832423, 56246211, 62117518, 148390399, 209085090, 10003248, 241313184, 25944135,
              212802310, 50222736, 18298478, 209886001, 145034471, 186841927, 160807241, 258257144,
              193915204, 92650808, 171362072, 30930936, 158727274, 226213489, 244216783, 158168844}))
  stage_3_butterfly_26 (
    .x_in(stage_2_per_out[52]),
    .y_in(stage_2_per_out[53]),
    .x_out(stage_3_per_in[52]),
    .y_out(stage_3_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({77981460, 199633043, 142181410, 160841949, 8411857, 100229847, 75073484, 13458851,
              192832423, 56246211, 62117518, 148390399, 209085090, 10003248, 241313184, 25944135,
              212802310, 50222736, 18298478, 209886001, 145034471, 186841927, 160807241, 258257144,
              193915204, 92650808, 171362072, 30930936, 158727274, 226213489, 244216783, 158168844}))
  stage_3_butterfly_27 (
    .x_in(stage_2_per_out[54]),
    .y_in(stage_2_per_out[55]),
    .x_out(stage_3_per_in[54]),
    .y_out(stage_3_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({77981460, 199633043, 142181410, 160841949, 8411857, 100229847, 75073484, 13458851,
              192832423, 56246211, 62117518, 148390399, 209085090, 10003248, 241313184, 25944135,
              212802310, 50222736, 18298478, 209886001, 145034471, 186841927, 160807241, 258257144,
              193915204, 92650808, 171362072, 30930936, 158727274, 226213489, 244216783, 158168844}))
  stage_3_butterfly_28 (
    .x_in(stage_2_per_out[56]),
    .y_in(stage_2_per_out[57]),
    .x_out(stage_3_per_in[56]),
    .y_out(stage_3_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({77981460, 199633043, 142181410, 160841949, 8411857, 100229847, 75073484, 13458851,
              192832423, 56246211, 62117518, 148390399, 209085090, 10003248, 241313184, 25944135,
              212802310, 50222736, 18298478, 209886001, 145034471, 186841927, 160807241, 258257144,
              193915204, 92650808, 171362072, 30930936, 158727274, 226213489, 244216783, 158168844}))
  stage_3_butterfly_29 (
    .x_in(stage_2_per_out[58]),
    .y_in(stage_2_per_out[59]),
    .x_out(stage_3_per_in[58]),
    .y_out(stage_3_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({77981460, 199633043, 142181410, 160841949, 8411857, 100229847, 75073484, 13458851,
              192832423, 56246211, 62117518, 148390399, 209085090, 10003248, 241313184, 25944135,
              212802310, 50222736, 18298478, 209886001, 145034471, 186841927, 160807241, 258257144,
              193915204, 92650808, 171362072, 30930936, 158727274, 226213489, 244216783, 158168844}))
  stage_3_butterfly_30 (
    .x_in(stage_2_per_out[60]),
    .y_in(stage_2_per_out[61]),
    .x_out(stage_3_per_in[60]),
    .y_out(stage_3_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({77981460, 199633043, 142181410, 160841949, 8411857, 100229847, 75073484, 13458851,
              192832423, 56246211, 62117518, 148390399, 209085090, 10003248, 241313184, 25944135,
              212802310, 50222736, 18298478, 209886001, 145034471, 186841927, 160807241, 258257144,
              193915204, 92650808, 171362072, 30930936, 158727274, 226213489, 244216783, 158168844}))
  stage_3_butterfly_31 (
    .x_in(stage_2_per_out[62]),
    .y_in(stage_2_per_out[63]),
    .x_out(stage_3_per_in[62]),
    .y_out(stage_3_per_in[63]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({219738759, 28242170, 132483080, 216395023, 42719459, 168676526, 212275822, 190319963,
              176209504, 138879618, 209725121, 66242139, 49057739, 262464837, 183029478, 80505160,
              202059197, 101414187, 200399539, 7460524, 34971158, 103234978, 206795535, 171051327,
              218231468, 143969870, 143779572, 211426643, 247253507, 242302870, 25853611, 36946189}))
  stage_3_butterfly_32 (
    .x_in(stage_2_per_out[64]),
    .y_in(stage_2_per_out[65]),
    .x_out(stage_3_per_in[64]),
    .y_out(stage_3_per_in[65]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({219738759, 28242170, 132483080, 216395023, 42719459, 168676526, 212275822, 190319963,
              176209504, 138879618, 209725121, 66242139, 49057739, 262464837, 183029478, 80505160,
              202059197, 101414187, 200399539, 7460524, 34971158, 103234978, 206795535, 171051327,
              218231468, 143969870, 143779572, 211426643, 247253507, 242302870, 25853611, 36946189}))
  stage_3_butterfly_33 (
    .x_in(stage_2_per_out[66]),
    .y_in(stage_2_per_out[67]),
    .x_out(stage_3_per_in[66]),
    .y_out(stage_3_per_in[67]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({219738759, 28242170, 132483080, 216395023, 42719459, 168676526, 212275822, 190319963,
              176209504, 138879618, 209725121, 66242139, 49057739, 262464837, 183029478, 80505160,
              202059197, 101414187, 200399539, 7460524, 34971158, 103234978, 206795535, 171051327,
              218231468, 143969870, 143779572, 211426643, 247253507, 242302870, 25853611, 36946189}))
  stage_3_butterfly_34 (
    .x_in(stage_2_per_out[68]),
    .y_in(stage_2_per_out[69]),
    .x_out(stage_3_per_in[68]),
    .y_out(stage_3_per_in[69]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({219738759, 28242170, 132483080, 216395023, 42719459, 168676526, 212275822, 190319963,
              176209504, 138879618, 209725121, 66242139, 49057739, 262464837, 183029478, 80505160,
              202059197, 101414187, 200399539, 7460524, 34971158, 103234978, 206795535, 171051327,
              218231468, 143969870, 143779572, 211426643, 247253507, 242302870, 25853611, 36946189}))
  stage_3_butterfly_35 (
    .x_in(stage_2_per_out[70]),
    .y_in(stage_2_per_out[71]),
    .x_out(stage_3_per_in[70]),
    .y_out(stage_3_per_in[71]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({219738759, 28242170, 132483080, 216395023, 42719459, 168676526, 212275822, 190319963,
              176209504, 138879618, 209725121, 66242139, 49057739, 262464837, 183029478, 80505160,
              202059197, 101414187, 200399539, 7460524, 34971158, 103234978, 206795535, 171051327,
              218231468, 143969870, 143779572, 211426643, 247253507, 242302870, 25853611, 36946189}))
  stage_3_butterfly_36 (
    .x_in(stage_2_per_out[72]),
    .y_in(stage_2_per_out[73]),
    .x_out(stage_3_per_in[72]),
    .y_out(stage_3_per_in[73]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({219738759, 28242170, 132483080, 216395023, 42719459, 168676526, 212275822, 190319963,
              176209504, 138879618, 209725121, 66242139, 49057739, 262464837, 183029478, 80505160,
              202059197, 101414187, 200399539, 7460524, 34971158, 103234978, 206795535, 171051327,
              218231468, 143969870, 143779572, 211426643, 247253507, 242302870, 25853611, 36946189}))
  stage_3_butterfly_37 (
    .x_in(stage_2_per_out[74]),
    .y_in(stage_2_per_out[75]),
    .x_out(stage_3_per_in[74]),
    .y_out(stage_3_per_in[75]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({219738759, 28242170, 132483080, 216395023, 42719459, 168676526, 212275822, 190319963,
              176209504, 138879618, 209725121, 66242139, 49057739, 262464837, 183029478, 80505160,
              202059197, 101414187, 200399539, 7460524, 34971158, 103234978, 206795535, 171051327,
              218231468, 143969870, 143779572, 211426643, 247253507, 242302870, 25853611, 36946189}))
  stage_3_butterfly_38 (
    .x_in(stage_2_per_out[76]),
    .y_in(stage_2_per_out[77]),
    .x_out(stage_3_per_in[76]),
    .y_out(stage_3_per_in[77]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({219738759, 28242170, 132483080, 216395023, 42719459, 168676526, 212275822, 190319963,
              176209504, 138879618, 209725121, 66242139, 49057739, 262464837, 183029478, 80505160,
              202059197, 101414187, 200399539, 7460524, 34971158, 103234978, 206795535, 171051327,
              218231468, 143969870, 143779572, 211426643, 247253507, 242302870, 25853611, 36946189}))
  stage_3_butterfly_39 (
    .x_in(stage_2_per_out[78]),
    .y_in(stage_2_per_out[79]),
    .x_out(stage_3_per_in[78]),
    .y_out(stage_3_per_in[79]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({24688427, 110403916, 170284131, 202071175, 224586596, 181281889, 205290416, 65413984,
              129576773, 61644903, 263077695, 67321994, 196771169, 82155735, 155060883, 207329882,
              258226806, 219898221, 167366585, 93469550, 68493159, 63483304, 225389748, 95251863,
              17231623, 252241817, 156366160, 35918322, 35924353, 6574921, 119169851, 6292910}))
  stage_3_butterfly_40 (
    .x_in(stage_2_per_out[80]),
    .y_in(stage_2_per_out[81]),
    .x_out(stage_3_per_in[80]),
    .y_out(stage_3_per_in[81]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({24688427, 110403916, 170284131, 202071175, 224586596, 181281889, 205290416, 65413984,
              129576773, 61644903, 263077695, 67321994, 196771169, 82155735, 155060883, 207329882,
              258226806, 219898221, 167366585, 93469550, 68493159, 63483304, 225389748, 95251863,
              17231623, 252241817, 156366160, 35918322, 35924353, 6574921, 119169851, 6292910}))
  stage_3_butterfly_41 (
    .x_in(stage_2_per_out[82]),
    .y_in(stage_2_per_out[83]),
    .x_out(stage_3_per_in[82]),
    .y_out(stage_3_per_in[83]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({24688427, 110403916, 170284131, 202071175, 224586596, 181281889, 205290416, 65413984,
              129576773, 61644903, 263077695, 67321994, 196771169, 82155735, 155060883, 207329882,
              258226806, 219898221, 167366585, 93469550, 68493159, 63483304, 225389748, 95251863,
              17231623, 252241817, 156366160, 35918322, 35924353, 6574921, 119169851, 6292910}))
  stage_3_butterfly_42 (
    .x_in(stage_2_per_out[84]),
    .y_in(stage_2_per_out[85]),
    .x_out(stage_3_per_in[84]),
    .y_out(stage_3_per_in[85]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({24688427, 110403916, 170284131, 202071175, 224586596, 181281889, 205290416, 65413984,
              129576773, 61644903, 263077695, 67321994, 196771169, 82155735, 155060883, 207329882,
              258226806, 219898221, 167366585, 93469550, 68493159, 63483304, 225389748, 95251863,
              17231623, 252241817, 156366160, 35918322, 35924353, 6574921, 119169851, 6292910}))
  stage_3_butterfly_43 (
    .x_in(stage_2_per_out[86]),
    .y_in(stage_2_per_out[87]),
    .x_out(stage_3_per_in[86]),
    .y_out(stage_3_per_in[87]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({24688427, 110403916, 170284131, 202071175, 224586596, 181281889, 205290416, 65413984,
              129576773, 61644903, 263077695, 67321994, 196771169, 82155735, 155060883, 207329882,
              258226806, 219898221, 167366585, 93469550, 68493159, 63483304, 225389748, 95251863,
              17231623, 252241817, 156366160, 35918322, 35924353, 6574921, 119169851, 6292910}))
  stage_3_butterfly_44 (
    .x_in(stage_2_per_out[88]),
    .y_in(stage_2_per_out[89]),
    .x_out(stage_3_per_in[88]),
    .y_out(stage_3_per_in[89]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({24688427, 110403916, 170284131, 202071175, 224586596, 181281889, 205290416, 65413984,
              129576773, 61644903, 263077695, 67321994, 196771169, 82155735, 155060883, 207329882,
              258226806, 219898221, 167366585, 93469550, 68493159, 63483304, 225389748, 95251863,
              17231623, 252241817, 156366160, 35918322, 35924353, 6574921, 119169851, 6292910}))
  stage_3_butterfly_45 (
    .x_in(stage_2_per_out[90]),
    .y_in(stage_2_per_out[91]),
    .x_out(stage_3_per_in[90]),
    .y_out(stage_3_per_in[91]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({24688427, 110403916, 170284131, 202071175, 224586596, 181281889, 205290416, 65413984,
              129576773, 61644903, 263077695, 67321994, 196771169, 82155735, 155060883, 207329882,
              258226806, 219898221, 167366585, 93469550, 68493159, 63483304, 225389748, 95251863,
              17231623, 252241817, 156366160, 35918322, 35924353, 6574921, 119169851, 6292910}))
  stage_3_butterfly_46 (
    .x_in(stage_2_per_out[92]),
    .y_in(stage_2_per_out[93]),
    .x_out(stage_3_per_in[92]),
    .y_out(stage_3_per_in[93]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({24688427, 110403916, 170284131, 202071175, 224586596, 181281889, 205290416, 65413984,
              129576773, 61644903, 263077695, 67321994, 196771169, 82155735, 155060883, 207329882,
              258226806, 219898221, 167366585, 93469550, 68493159, 63483304, 225389748, 95251863,
              17231623, 252241817, 156366160, 35918322, 35924353, 6574921, 119169851, 6292910}))
  stage_3_butterfly_47 (
    .x_in(stage_2_per_out[94]),
    .y_in(stage_2_per_out[95]),
    .x_out(stage_3_per_in[94]),
    .y_out(stage_3_per_in[95]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({4839268, 178386996, 102915173, 167911982, 263070789, 131377029, 82934386, 76925614,
              117274103, 73081523, 68267735, 68559335, 55609416, 190980049, 243024363, 195748297,
              10720790, 210770212, 236109059, 222861227, 225265815, 256272276, 47879495, 177340471,
              40718170, 165350229, 43194148, 200749611, 256869432, 209583375, 139268485, 257269778}))
  stage_3_butterfly_48 (
    .x_in(stage_2_per_out[96]),
    .y_in(stage_2_per_out[97]),
    .x_out(stage_3_per_in[96]),
    .y_out(stage_3_per_in[97]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({4839268, 178386996, 102915173, 167911982, 263070789, 131377029, 82934386, 76925614,
              117274103, 73081523, 68267735, 68559335, 55609416, 190980049, 243024363, 195748297,
              10720790, 210770212, 236109059, 222861227, 225265815, 256272276, 47879495, 177340471,
              40718170, 165350229, 43194148, 200749611, 256869432, 209583375, 139268485, 257269778}))
  stage_3_butterfly_49 (
    .x_in(stage_2_per_out[98]),
    .y_in(stage_2_per_out[99]),
    .x_out(stage_3_per_in[98]),
    .y_out(stage_3_per_in[99]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({4839268, 178386996, 102915173, 167911982, 263070789, 131377029, 82934386, 76925614,
              117274103, 73081523, 68267735, 68559335, 55609416, 190980049, 243024363, 195748297,
              10720790, 210770212, 236109059, 222861227, 225265815, 256272276, 47879495, 177340471,
              40718170, 165350229, 43194148, 200749611, 256869432, 209583375, 139268485, 257269778}))
  stage_3_butterfly_50 (
    .x_in(stage_2_per_out[100]),
    .y_in(stage_2_per_out[101]),
    .x_out(stage_3_per_in[100]),
    .y_out(stage_3_per_in[101]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({4839268, 178386996, 102915173, 167911982, 263070789, 131377029, 82934386, 76925614,
              117274103, 73081523, 68267735, 68559335, 55609416, 190980049, 243024363, 195748297,
              10720790, 210770212, 236109059, 222861227, 225265815, 256272276, 47879495, 177340471,
              40718170, 165350229, 43194148, 200749611, 256869432, 209583375, 139268485, 257269778}))
  stage_3_butterfly_51 (
    .x_in(stage_2_per_out[102]),
    .y_in(stage_2_per_out[103]),
    .x_out(stage_3_per_in[102]),
    .y_out(stage_3_per_in[103]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({4839268, 178386996, 102915173, 167911982, 263070789, 131377029, 82934386, 76925614,
              117274103, 73081523, 68267735, 68559335, 55609416, 190980049, 243024363, 195748297,
              10720790, 210770212, 236109059, 222861227, 225265815, 256272276, 47879495, 177340471,
              40718170, 165350229, 43194148, 200749611, 256869432, 209583375, 139268485, 257269778}))
  stage_3_butterfly_52 (
    .x_in(stage_2_per_out[104]),
    .y_in(stage_2_per_out[105]),
    .x_out(stage_3_per_in[104]),
    .y_out(stage_3_per_in[105]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({4839268, 178386996, 102915173, 167911982, 263070789, 131377029, 82934386, 76925614,
              117274103, 73081523, 68267735, 68559335, 55609416, 190980049, 243024363, 195748297,
              10720790, 210770212, 236109059, 222861227, 225265815, 256272276, 47879495, 177340471,
              40718170, 165350229, 43194148, 200749611, 256869432, 209583375, 139268485, 257269778}))
  stage_3_butterfly_53 (
    .x_in(stage_2_per_out[106]),
    .y_in(stage_2_per_out[107]),
    .x_out(stage_3_per_in[106]),
    .y_out(stage_3_per_in[107]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({4839268, 178386996, 102915173, 167911982, 263070789, 131377029, 82934386, 76925614,
              117274103, 73081523, 68267735, 68559335, 55609416, 190980049, 243024363, 195748297,
              10720790, 210770212, 236109059, 222861227, 225265815, 256272276, 47879495, 177340471,
              40718170, 165350229, 43194148, 200749611, 256869432, 209583375, 139268485, 257269778}))
  stage_3_butterfly_54 (
    .x_in(stage_2_per_out[108]),
    .y_in(stage_2_per_out[109]),
    .x_out(stage_3_per_in[108]),
    .y_out(stage_3_per_in[109]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({4839268, 178386996, 102915173, 167911982, 263070789, 131377029, 82934386, 76925614,
              117274103, 73081523, 68267735, 68559335, 55609416, 190980049, 243024363, 195748297,
              10720790, 210770212, 236109059, 222861227, 225265815, 256272276, 47879495, 177340471,
              40718170, 165350229, 43194148, 200749611, 256869432, 209583375, 139268485, 257269778}))
  stage_3_butterfly_55 (
    .x_in(stage_2_per_out[110]),
    .y_in(stage_2_per_out[111]),
    .x_out(stage_3_per_in[110]),
    .y_out(stage_3_per_in[111]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({233888407, 23405380, 169182486, 254132077, 34256894, 79136411, 109479656, 205525433,
              60548134, 140366124, 210734246, 149992379, 50986641, 114486793, 266671862, 184310992,
              237102043, 131023241, 229100654, 196522490, 185138250, 122332647, 247289727, 196328787,
              154421517, 238382196, 171541778, 61997323, 242025902, 137672988, 49675259, 182691070}))
  stage_3_butterfly_56 (
    .x_in(stage_2_per_out[112]),
    .y_in(stage_2_per_out[113]),
    .x_out(stage_3_per_in[112]),
    .y_out(stage_3_per_in[113]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({233888407, 23405380, 169182486, 254132077, 34256894, 79136411, 109479656, 205525433,
              60548134, 140366124, 210734246, 149992379, 50986641, 114486793, 266671862, 184310992,
              237102043, 131023241, 229100654, 196522490, 185138250, 122332647, 247289727, 196328787,
              154421517, 238382196, 171541778, 61997323, 242025902, 137672988, 49675259, 182691070}))
  stage_3_butterfly_57 (
    .x_in(stage_2_per_out[114]),
    .y_in(stage_2_per_out[115]),
    .x_out(stage_3_per_in[114]),
    .y_out(stage_3_per_in[115]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({233888407, 23405380, 169182486, 254132077, 34256894, 79136411, 109479656, 205525433,
              60548134, 140366124, 210734246, 149992379, 50986641, 114486793, 266671862, 184310992,
              237102043, 131023241, 229100654, 196522490, 185138250, 122332647, 247289727, 196328787,
              154421517, 238382196, 171541778, 61997323, 242025902, 137672988, 49675259, 182691070}))
  stage_3_butterfly_58 (
    .x_in(stage_2_per_out[116]),
    .y_in(stage_2_per_out[117]),
    .x_out(stage_3_per_in[116]),
    .y_out(stage_3_per_in[117]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({233888407, 23405380, 169182486, 254132077, 34256894, 79136411, 109479656, 205525433,
              60548134, 140366124, 210734246, 149992379, 50986641, 114486793, 266671862, 184310992,
              237102043, 131023241, 229100654, 196522490, 185138250, 122332647, 247289727, 196328787,
              154421517, 238382196, 171541778, 61997323, 242025902, 137672988, 49675259, 182691070}))
  stage_3_butterfly_59 (
    .x_in(stage_2_per_out[118]),
    .y_in(stage_2_per_out[119]),
    .x_out(stage_3_per_in[118]),
    .y_out(stage_3_per_in[119]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({233888407, 23405380, 169182486, 254132077, 34256894, 79136411, 109479656, 205525433,
              60548134, 140366124, 210734246, 149992379, 50986641, 114486793, 266671862, 184310992,
              237102043, 131023241, 229100654, 196522490, 185138250, 122332647, 247289727, 196328787,
              154421517, 238382196, 171541778, 61997323, 242025902, 137672988, 49675259, 182691070}))
  stage_3_butterfly_60 (
    .x_in(stage_2_per_out[120]),
    .y_in(stage_2_per_out[121]),
    .x_out(stage_3_per_in[120]),
    .y_out(stage_3_per_in[121]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({233888407, 23405380, 169182486, 254132077, 34256894, 79136411, 109479656, 205525433,
              60548134, 140366124, 210734246, 149992379, 50986641, 114486793, 266671862, 184310992,
              237102043, 131023241, 229100654, 196522490, 185138250, 122332647, 247289727, 196328787,
              154421517, 238382196, 171541778, 61997323, 242025902, 137672988, 49675259, 182691070}))
  stage_3_butterfly_61 (
    .x_in(stage_2_per_out[122]),
    .y_in(stage_2_per_out[123]),
    .x_out(stage_3_per_in[122]),
    .y_out(stage_3_per_in[123]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({233888407, 23405380, 169182486, 254132077, 34256894, 79136411, 109479656, 205525433,
              60548134, 140366124, 210734246, 149992379, 50986641, 114486793, 266671862, 184310992,
              237102043, 131023241, 229100654, 196522490, 185138250, 122332647, 247289727, 196328787,
              154421517, 238382196, 171541778, 61997323, 242025902, 137672988, 49675259, 182691070}))
  stage_3_butterfly_62 (
    .x_in(stage_2_per_out[124]),
    .y_in(stage_2_per_out[125]),
    .x_out(stage_3_per_in[124]),
    .y_out(stage_3_per_in[125]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({233888407, 23405380, 169182486, 254132077, 34256894, 79136411, 109479656, 205525433,
              60548134, 140366124, 210734246, 149992379, 50986641, 114486793, 266671862, 184310992,
              237102043, 131023241, 229100654, 196522490, 185138250, 122332647, 247289727, 196328787,
              154421517, 238382196, 171541778, 61997323, 242025902, 137672988, 49675259, 182691070}))
  stage_3_butterfly_63 (
    .x_in(stage_2_per_out[126]),
    .y_in(stage_2_per_out[127]),
    .x_out(stage_3_per_in[126]),
    .y_out(stage_3_per_in[127]),
    .clk(clk),
    .rst(rst)
  );



  // TODO(Yang): stage 3 -> stage 4 permutation
  // FIXME: ignore butterfly units for now.
  stage_3_permutation #(
    .DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    .INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_3_4_per (
    .inData_0(stage_3_per_in[0]),
    .inData_1(stage_3_per_in[1]),
    .inData_2(stage_3_per_in[2]),
    .inData_3(stage_3_per_in[3]),
    .inData_4(stage_3_per_in[4]),
    .inData_5(stage_3_per_in[5]),
    .inData_6(stage_3_per_in[6]),
    .inData_7(stage_3_per_in[7]),
    .inData_8(stage_3_per_in[8]),
    .inData_9(stage_3_per_in[9]),
    .inData_10(stage_3_per_in[10]),
    .inData_11(stage_3_per_in[11]),
    .inData_12(stage_3_per_in[12]),
    .inData_13(stage_3_per_in[13]),
    .inData_14(stage_3_per_in[14]),
    .inData_15(stage_3_per_in[15]),
    .inData_16(stage_3_per_in[16]),
    .inData_17(stage_3_per_in[17]),
    .inData_18(stage_3_per_in[18]),
    .inData_19(stage_3_per_in[19]),
    .inData_20(stage_3_per_in[20]),
    .inData_21(stage_3_per_in[21]),
    .inData_22(stage_3_per_in[22]),
    .inData_23(stage_3_per_in[23]),
    .inData_24(stage_3_per_in[24]),
    .inData_25(stage_3_per_in[25]),
    .inData_26(stage_3_per_in[26]),
    .inData_27(stage_3_per_in[27]),
    .inData_28(stage_3_per_in[28]),
    .inData_29(stage_3_per_in[29]),
    .inData_30(stage_3_per_in[30]),
    .inData_31(stage_3_per_in[31]),
    .inData_32(stage_3_per_in[32]),
    .inData_33(stage_3_per_in[33]),
    .inData_34(stage_3_per_in[34]),
    .inData_35(stage_3_per_in[35]),
    .inData_36(stage_3_per_in[36]),
    .inData_37(stage_3_per_in[37]),
    .inData_38(stage_3_per_in[38]),
    .inData_39(stage_3_per_in[39]),
    .inData_40(stage_3_per_in[40]),
    .inData_41(stage_3_per_in[41]),
    .inData_42(stage_3_per_in[42]),
    .inData_43(stage_3_per_in[43]),
    .inData_44(stage_3_per_in[44]),
    .inData_45(stage_3_per_in[45]),
    .inData_46(stage_3_per_in[46]),
    .inData_47(stage_3_per_in[47]),
    .inData_48(stage_3_per_in[48]),
    .inData_49(stage_3_per_in[49]),
    .inData_50(stage_3_per_in[50]),
    .inData_51(stage_3_per_in[51]),
    .inData_52(stage_3_per_in[52]),
    .inData_53(stage_3_per_in[53]),
    .inData_54(stage_3_per_in[54]),
    .inData_55(stage_3_per_in[55]),
    .inData_56(stage_3_per_in[56]),
    .inData_57(stage_3_per_in[57]),
    .inData_58(stage_3_per_in[58]),
    .inData_59(stage_3_per_in[59]),
    .inData_60(stage_3_per_in[60]),
    .inData_61(stage_3_per_in[61]),
    .inData_62(stage_3_per_in[62]),
    .inData_63(stage_3_per_in[63]),
    .inData_64(stage_3_per_in[64]),
    .inData_65(stage_3_per_in[65]),
    .inData_66(stage_3_per_in[66]),
    .inData_67(stage_3_per_in[67]),
    .inData_68(stage_3_per_in[68]),
    .inData_69(stage_3_per_in[69]),
    .inData_70(stage_3_per_in[70]),
    .inData_71(stage_3_per_in[71]),
    .inData_72(stage_3_per_in[72]),
    .inData_73(stage_3_per_in[73]),
    .inData_74(stage_3_per_in[74]),
    .inData_75(stage_3_per_in[75]),
    .inData_76(stage_3_per_in[76]),
    .inData_77(stage_3_per_in[77]),
    .inData_78(stage_3_per_in[78]),
    .inData_79(stage_3_per_in[79]),
    .inData_80(stage_3_per_in[80]),
    .inData_81(stage_3_per_in[81]),
    .inData_82(stage_3_per_in[82]),
    .inData_83(stage_3_per_in[83]),
    .inData_84(stage_3_per_in[84]),
    .inData_85(stage_3_per_in[85]),
    .inData_86(stage_3_per_in[86]),
    .inData_87(stage_3_per_in[87]),
    .inData_88(stage_3_per_in[88]),
    .inData_89(stage_3_per_in[89]),
    .inData_90(stage_3_per_in[90]),
    .inData_91(stage_3_per_in[91]),
    .inData_92(stage_3_per_in[92]),
    .inData_93(stage_3_per_in[93]),
    .inData_94(stage_3_per_in[94]),
    .inData_95(stage_3_per_in[95]),
    .inData_96(stage_3_per_in[96]),
    .inData_97(stage_3_per_in[97]),
    .inData_98(stage_3_per_in[98]),
    .inData_99(stage_3_per_in[99]),
    .inData_100(stage_3_per_in[100]),
    .inData_101(stage_3_per_in[101]),
    .inData_102(stage_3_per_in[102]),
    .inData_103(stage_3_per_in[103]),
    .inData_104(stage_3_per_in[104]),
    .inData_105(stage_3_per_in[105]),
    .inData_106(stage_3_per_in[106]),
    .inData_107(stage_3_per_in[107]),
    .inData_108(stage_3_per_in[108]),
    .inData_109(stage_3_per_in[109]),
    .inData_110(stage_3_per_in[110]),
    .inData_111(stage_3_per_in[111]),
    .inData_112(stage_3_per_in[112]),
    .inData_113(stage_3_per_in[113]),
    .inData_114(stage_3_per_in[114]),
    .inData_115(stage_3_per_in[115]),
    .inData_116(stage_3_per_in[116]),
    .inData_117(stage_3_per_in[117]),
    .inData_118(stage_3_per_in[118]),
    .inData_119(stage_3_per_in[119]),
    .inData_120(stage_3_per_in[120]),
    .inData_121(stage_3_per_in[121]),
    .inData_122(stage_3_per_in[122]),
    .inData_123(stage_3_per_in[123]),
    .inData_124(stage_3_per_in[124]),
    .inData_125(stage_3_per_in[125]),
    .inData_126(stage_3_per_in[126]),
    .inData_127(stage_3_per_in[127]),
    .outData_0(stage_3_per_out[0]),
    .outData_1(stage_3_per_out[1]),
    .outData_2(stage_3_per_out[2]),
    .outData_3(stage_3_per_out[3]),
    .outData_4(stage_3_per_out[4]),
    .outData_5(stage_3_per_out[5]),
    .outData_6(stage_3_per_out[6]),
    .outData_7(stage_3_per_out[7]),
    .outData_8(stage_3_per_out[8]),
    .outData_9(stage_3_per_out[9]),
    .outData_10(stage_3_per_out[10]),
    .outData_11(stage_3_per_out[11]),
    .outData_12(stage_3_per_out[12]),
    .outData_13(stage_3_per_out[13]),
    .outData_14(stage_3_per_out[14]),
    .outData_15(stage_3_per_out[15]),
    .outData_16(stage_3_per_out[16]),
    .outData_17(stage_3_per_out[17]),
    .outData_18(stage_3_per_out[18]),
    .outData_19(stage_3_per_out[19]),
    .outData_20(stage_3_per_out[20]),
    .outData_21(stage_3_per_out[21]),
    .outData_22(stage_3_per_out[22]),
    .outData_23(stage_3_per_out[23]),
    .outData_24(stage_3_per_out[24]),
    .outData_25(stage_3_per_out[25]),
    .outData_26(stage_3_per_out[26]),
    .outData_27(stage_3_per_out[27]),
    .outData_28(stage_3_per_out[28]),
    .outData_29(stage_3_per_out[29]),
    .outData_30(stage_3_per_out[30]),
    .outData_31(stage_3_per_out[31]),
    .outData_32(stage_3_per_out[32]),
    .outData_33(stage_3_per_out[33]),
    .outData_34(stage_3_per_out[34]),
    .outData_35(stage_3_per_out[35]),
    .outData_36(stage_3_per_out[36]),
    .outData_37(stage_3_per_out[37]),
    .outData_38(stage_3_per_out[38]),
    .outData_39(stage_3_per_out[39]),
    .outData_40(stage_3_per_out[40]),
    .outData_41(stage_3_per_out[41]),
    .outData_42(stage_3_per_out[42]),
    .outData_43(stage_3_per_out[43]),
    .outData_44(stage_3_per_out[44]),
    .outData_45(stage_3_per_out[45]),
    .outData_46(stage_3_per_out[46]),
    .outData_47(stage_3_per_out[47]),
    .outData_48(stage_3_per_out[48]),
    .outData_49(stage_3_per_out[49]),
    .outData_50(stage_3_per_out[50]),
    .outData_51(stage_3_per_out[51]),
    .outData_52(stage_3_per_out[52]),
    .outData_53(stage_3_per_out[53]),
    .outData_54(stage_3_per_out[54]),
    .outData_55(stage_3_per_out[55]),
    .outData_56(stage_3_per_out[56]),
    .outData_57(stage_3_per_out[57]),
    .outData_58(stage_3_per_out[58]),
    .outData_59(stage_3_per_out[59]),
    .outData_60(stage_3_per_out[60]),
    .outData_61(stage_3_per_out[61]),
    .outData_62(stage_3_per_out[62]),
    .outData_63(stage_3_per_out[63]),
    .outData_64(stage_3_per_out[64]),
    .outData_65(stage_3_per_out[65]),
    .outData_66(stage_3_per_out[66]),
    .outData_67(stage_3_per_out[67]),
    .outData_68(stage_3_per_out[68]),
    .outData_69(stage_3_per_out[69]),
    .outData_70(stage_3_per_out[70]),
    .outData_71(stage_3_per_out[71]),
    .outData_72(stage_3_per_out[72]),
    .outData_73(stage_3_per_out[73]),
    .outData_74(stage_3_per_out[74]),
    .outData_75(stage_3_per_out[75]),
    .outData_76(stage_3_per_out[76]),
    .outData_77(stage_3_per_out[77]),
    .outData_78(stage_3_per_out[78]),
    .outData_79(stage_3_per_out[79]),
    .outData_80(stage_3_per_out[80]),
    .outData_81(stage_3_per_out[81]),
    .outData_82(stage_3_per_out[82]),
    .outData_83(stage_3_per_out[83]),
    .outData_84(stage_3_per_out[84]),
    .outData_85(stage_3_per_out[85]),
    .outData_86(stage_3_per_out[86]),
    .outData_87(stage_3_per_out[87]),
    .outData_88(stage_3_per_out[88]),
    .outData_89(stage_3_per_out[89]),
    .outData_90(stage_3_per_out[90]),
    .outData_91(stage_3_per_out[91]),
    .outData_92(stage_3_per_out[92]),
    .outData_93(stage_3_per_out[93]),
    .outData_94(stage_3_per_out[94]),
    .outData_95(stage_3_per_out[95]),
    .outData_96(stage_3_per_out[96]),
    .outData_97(stage_3_per_out[97]),
    .outData_98(stage_3_per_out[98]),
    .outData_99(stage_3_per_out[99]),
    .outData_100(stage_3_per_out[100]),
    .outData_101(stage_3_per_out[101]),
    .outData_102(stage_3_per_out[102]),
    .outData_103(stage_3_per_out[103]),
    .outData_104(stage_3_per_out[104]),
    .outData_105(stage_3_per_out[105]),
    .outData_106(stage_3_per_out[106]),
    .outData_107(stage_3_per_out[107]),
    .outData_108(stage_3_per_out[108]),
    .outData_109(stage_3_per_out[109]),
    .outData_110(stage_3_per_out[110]),
    .outData_111(stage_3_per_out[111]),
    .outData_112(stage_3_per_out[112]),
    .outData_113(stage_3_per_out[113]),
    .outData_114(stage_3_per_out[114]),
    .outData_115(stage_3_per_out[115]),
    .outData_116(stage_3_per_out[116]),
    .outData_117(stage_3_per_out[117]),
    .outData_118(stage_3_per_out[118]),
    .outData_119(stage_3_per_out[119]),
    .outData_120(stage_3_per_out[120]),
    .outData_121(stage_3_per_out[121]),
    .outData_122(stage_3_per_out[122]),
    .outData_123(stage_3_per_out[123]),
    .outData_124(stage_3_per_out[124]),
    .outData_125(stage_3_per_out[125]),
    .outData_126(stage_3_per_out[126]),
    .outData_127(stage_3_per_out[127]),
    .in_start(in_start[3]),
    .out_start(out_start[3]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 4 32 butterfly units
  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 11101448, 189762285, 244883276, 229228230, 101839787, 85922744, 10571783,
              117496916, 192696288, 106640438, 90597117, 189881206, 241125460, 209161759, 245906264,
              55721255, 64217206, 40553702, 214551729, 226739459, 246744565, 104557084, 104784816,
              122008382, 225636920, 47994339, 168407516, 184226747, 69161747, 239545014, 72738487}))
  stage_4_butterfly_0 (
    .x_in(stage_3_per_out[0]),
    .y_in(stage_3_per_out[1]),
    .x_out(stage_4_per_in[0]),
    .y_out(stage_4_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 11101448, 189762285, 244883276, 229228230, 101839787, 85922744, 10571783,
              117496916, 192696288, 106640438, 90597117, 189881206, 241125460, 209161759, 245906264,
              55721255, 64217206, 40553702, 214551729, 226739459, 246744565, 104557084, 104784816,
              122008382, 225636920, 47994339, 168407516, 184226747, 69161747, 239545014, 72738487}))
  stage_4_butterfly_1 (
    .x_in(stage_3_per_out[2]),
    .y_in(stage_3_per_out[3]),
    .x_out(stage_4_per_in[2]),
    .y_out(stage_4_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 11101448, 189762285, 244883276, 229228230, 101839787, 85922744, 10571783,
              117496916, 192696288, 106640438, 90597117, 189881206, 241125460, 209161759, 245906264,
              55721255, 64217206, 40553702, 214551729, 226739459, 246744565, 104557084, 104784816,
              122008382, 225636920, 47994339, 168407516, 184226747, 69161747, 239545014, 72738487}))
  stage_4_butterfly_2 (
    .x_in(stage_3_per_out[4]),
    .y_in(stage_3_per_out[5]),
    .x_out(stage_4_per_in[4]),
    .y_out(stage_4_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 11101448, 189762285, 244883276, 229228230, 101839787, 85922744, 10571783,
              117496916, 192696288, 106640438, 90597117, 189881206, 241125460, 209161759, 245906264,
              55721255, 64217206, 40553702, 214551729, 226739459, 246744565, 104557084, 104784816,
              122008382, 225636920, 47994339, 168407516, 184226747, 69161747, 239545014, 72738487}))
  stage_4_butterfly_3 (
    .x_in(stage_3_per_out[6]),
    .y_in(stage_3_per_out[7]),
    .x_out(stage_4_per_in[6]),
    .y_out(stage_4_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 11101448, 189762285, 244883276, 229228230, 101839787, 85922744, 10571783,
              117496916, 192696288, 106640438, 90597117, 189881206, 241125460, 209161759, 245906264,
              55721255, 64217206, 40553702, 214551729, 226739459, 246744565, 104557084, 104784816,
              122008382, 225636920, 47994339, 168407516, 184226747, 69161747, 239545014, 72738487}))
  stage_4_butterfly_4 (
    .x_in(stage_3_per_out[8]),
    .y_in(stage_3_per_out[9]),
    .x_out(stage_4_per_in[8]),
    .y_out(stage_4_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 11101448, 189762285, 244883276, 229228230, 101839787, 85922744, 10571783,
              117496916, 192696288, 106640438, 90597117, 189881206, 241125460, 209161759, 245906264,
              55721255, 64217206, 40553702, 214551729, 226739459, 246744565, 104557084, 104784816,
              122008382, 225636920, 47994339, 168407516, 184226747, 69161747, 239545014, 72738487}))
  stage_4_butterfly_5 (
    .x_in(stage_3_per_out[10]),
    .y_in(stage_3_per_out[11]),
    .x_out(stage_4_per_in[10]),
    .y_out(stage_4_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 11101448, 189762285, 244883276, 229228230, 101839787, 85922744, 10571783,
              117496916, 192696288, 106640438, 90597117, 189881206, 241125460, 209161759, 245906264,
              55721255, 64217206, 40553702, 214551729, 226739459, 246744565, 104557084, 104784816,
              122008382, 225636920, 47994339, 168407516, 184226747, 69161747, 239545014, 72738487}))
  stage_4_butterfly_6 (
    .x_in(stage_3_per_out[12]),
    .y_in(stage_3_per_out[13]),
    .x_out(stage_4_per_in[12]),
    .y_out(stage_4_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 11101448, 189762285, 244883276, 229228230, 101839787, 85922744, 10571783,
              117496916, 192696288, 106640438, 90597117, 189881206, 241125460, 209161759, 245906264,
              55721255, 64217206, 40553702, 214551729, 226739459, 246744565, 104557084, 104784816,
              122008382, 225636920, 47994339, 168407516, 184226747, 69161747, 239545014, 72738487}))
  stage_4_butterfly_7 (
    .x_in(stage_3_per_out[14]),
    .y_in(stage_3_per_out[15]),
    .x_out(stage_4_per_in[14]),
    .y_out(stage_4_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 11101448, 189762285, 244883276, 229228230, 101839787, 85922744, 10571783,
              117496916, 192696288, 106640438, 90597117, 189881206, 241125460, 209161759, 245906264,
              55721255, 64217206, 40553702, 214551729, 226739459, 246744565, 104557084, 104784816,
              122008382, 225636920, 47994339, 168407516, 184226747, 69161747, 239545014, 72738487}))
  stage_4_butterfly_8 (
    .x_in(stage_3_per_out[16]),
    .y_in(stage_3_per_out[17]),
    .x_out(stage_4_per_in[16]),
    .y_out(stage_4_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 11101448, 189762285, 244883276, 229228230, 101839787, 85922744, 10571783,
              117496916, 192696288, 106640438, 90597117, 189881206, 241125460, 209161759, 245906264,
              55721255, 64217206, 40553702, 214551729, 226739459, 246744565, 104557084, 104784816,
              122008382, 225636920, 47994339, 168407516, 184226747, 69161747, 239545014, 72738487}))
  stage_4_butterfly_9 (
    .x_in(stage_3_per_out[18]),
    .y_in(stage_3_per_out[19]),
    .x_out(stage_4_per_in[18]),
    .y_out(stage_4_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 11101448, 189762285, 244883276, 229228230, 101839787, 85922744, 10571783,
              117496916, 192696288, 106640438, 90597117, 189881206, 241125460, 209161759, 245906264,
              55721255, 64217206, 40553702, 214551729, 226739459, 246744565, 104557084, 104784816,
              122008382, 225636920, 47994339, 168407516, 184226747, 69161747, 239545014, 72738487}))
  stage_4_butterfly_10 (
    .x_in(stage_3_per_out[20]),
    .y_in(stage_3_per_out[21]),
    .x_out(stage_4_per_in[20]),
    .y_out(stage_4_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 11101448, 189762285, 244883276, 229228230, 101839787, 85922744, 10571783,
              117496916, 192696288, 106640438, 90597117, 189881206, 241125460, 209161759, 245906264,
              55721255, 64217206, 40553702, 214551729, 226739459, 246744565, 104557084, 104784816,
              122008382, 225636920, 47994339, 168407516, 184226747, 69161747, 239545014, 72738487}))
  stage_4_butterfly_11 (
    .x_in(stage_3_per_out[22]),
    .y_in(stage_3_per_out[23]),
    .x_out(stage_4_per_in[22]),
    .y_out(stage_4_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 11101448, 189762285, 244883276, 229228230, 101839787, 85922744, 10571783,
              117496916, 192696288, 106640438, 90597117, 189881206, 241125460, 209161759, 245906264,
              55721255, 64217206, 40553702, 214551729, 226739459, 246744565, 104557084, 104784816,
              122008382, 225636920, 47994339, 168407516, 184226747, 69161747, 239545014, 72738487}))
  stage_4_butterfly_12 (
    .x_in(stage_3_per_out[24]),
    .y_in(stage_3_per_out[25]),
    .x_out(stage_4_per_in[24]),
    .y_out(stage_4_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 11101448, 189762285, 244883276, 229228230, 101839787, 85922744, 10571783,
              117496916, 192696288, 106640438, 90597117, 189881206, 241125460, 209161759, 245906264,
              55721255, 64217206, 40553702, 214551729, 226739459, 246744565, 104557084, 104784816,
              122008382, 225636920, 47994339, 168407516, 184226747, 69161747, 239545014, 72738487}))
  stage_4_butterfly_13 (
    .x_in(stage_3_per_out[26]),
    .y_in(stage_3_per_out[27]),
    .x_out(stage_4_per_in[26]),
    .y_out(stage_4_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 11101448, 189762285, 244883276, 229228230, 101839787, 85922744, 10571783,
              117496916, 192696288, 106640438, 90597117, 189881206, 241125460, 209161759, 245906264,
              55721255, 64217206, 40553702, 214551729, 226739459, 246744565, 104557084, 104784816,
              122008382, 225636920, 47994339, 168407516, 184226747, 69161747, 239545014, 72738487}))
  stage_4_butterfly_14 (
    .x_in(stage_3_per_out[28]),
    .y_in(stage_3_per_out[29]),
    .x_out(stage_4_per_in[28]),
    .y_out(stage_4_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 11101448, 189762285, 244883276, 229228230, 101839787, 85922744, 10571783,
              117496916, 192696288, 106640438, 90597117, 189881206, 241125460, 209161759, 245906264,
              55721255, 64217206, 40553702, 214551729, 226739459, 246744565, 104557084, 104784816,
              122008382, 225636920, 47994339, 168407516, 184226747, 69161747, 239545014, 72738487}))
  stage_4_butterfly_15 (
    .x_in(stage_3_per_out[30]),
    .y_in(stage_3_per_out[31]),
    .x_out(stage_4_per_in[30]),
    .y_out(stage_4_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 68136911, 21713495, 7055647, 148662095, 256040960, 123185272, 170227406,
              193371292, 159404461, 183348420, 173702965, 186592442, 243304319, 236144340, 189591954,
              254509489, 66148505, 118518376, 108810259, 67012048, 104174682, 155168409, 3883583,
              25569479, 120936039, 13519489, 132703565, 71933862, 180525688, 139555205, 171721518}))
  stage_4_butterfly_16 (
    .x_in(stage_3_per_out[32]),
    .y_in(stage_3_per_out[33]),
    .x_out(stage_4_per_in[32]),
    .y_out(stage_4_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 68136911, 21713495, 7055647, 148662095, 256040960, 123185272, 170227406,
              193371292, 159404461, 183348420, 173702965, 186592442, 243304319, 236144340, 189591954,
              254509489, 66148505, 118518376, 108810259, 67012048, 104174682, 155168409, 3883583,
              25569479, 120936039, 13519489, 132703565, 71933862, 180525688, 139555205, 171721518}))
  stage_4_butterfly_17 (
    .x_in(stage_3_per_out[34]),
    .y_in(stage_3_per_out[35]),
    .x_out(stage_4_per_in[34]),
    .y_out(stage_4_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 68136911, 21713495, 7055647, 148662095, 256040960, 123185272, 170227406,
              193371292, 159404461, 183348420, 173702965, 186592442, 243304319, 236144340, 189591954,
              254509489, 66148505, 118518376, 108810259, 67012048, 104174682, 155168409, 3883583,
              25569479, 120936039, 13519489, 132703565, 71933862, 180525688, 139555205, 171721518}))
  stage_4_butterfly_18 (
    .x_in(stage_3_per_out[36]),
    .y_in(stage_3_per_out[37]),
    .x_out(stage_4_per_in[36]),
    .y_out(stage_4_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 68136911, 21713495, 7055647, 148662095, 256040960, 123185272, 170227406,
              193371292, 159404461, 183348420, 173702965, 186592442, 243304319, 236144340, 189591954,
              254509489, 66148505, 118518376, 108810259, 67012048, 104174682, 155168409, 3883583,
              25569479, 120936039, 13519489, 132703565, 71933862, 180525688, 139555205, 171721518}))
  stage_4_butterfly_19 (
    .x_in(stage_3_per_out[38]),
    .y_in(stage_3_per_out[39]),
    .x_out(stage_4_per_in[38]),
    .y_out(stage_4_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 68136911, 21713495, 7055647, 148662095, 256040960, 123185272, 170227406,
              193371292, 159404461, 183348420, 173702965, 186592442, 243304319, 236144340, 189591954,
              254509489, 66148505, 118518376, 108810259, 67012048, 104174682, 155168409, 3883583,
              25569479, 120936039, 13519489, 132703565, 71933862, 180525688, 139555205, 171721518}))
  stage_4_butterfly_20 (
    .x_in(stage_3_per_out[40]),
    .y_in(stage_3_per_out[41]),
    .x_out(stage_4_per_in[40]),
    .y_out(stage_4_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 68136911, 21713495, 7055647, 148662095, 256040960, 123185272, 170227406,
              193371292, 159404461, 183348420, 173702965, 186592442, 243304319, 236144340, 189591954,
              254509489, 66148505, 118518376, 108810259, 67012048, 104174682, 155168409, 3883583,
              25569479, 120936039, 13519489, 132703565, 71933862, 180525688, 139555205, 171721518}))
  stage_4_butterfly_21 (
    .x_in(stage_3_per_out[42]),
    .y_in(stage_3_per_out[43]),
    .x_out(stage_4_per_in[42]),
    .y_out(stage_4_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 68136911, 21713495, 7055647, 148662095, 256040960, 123185272, 170227406,
              193371292, 159404461, 183348420, 173702965, 186592442, 243304319, 236144340, 189591954,
              254509489, 66148505, 118518376, 108810259, 67012048, 104174682, 155168409, 3883583,
              25569479, 120936039, 13519489, 132703565, 71933862, 180525688, 139555205, 171721518}))
  stage_4_butterfly_22 (
    .x_in(stage_3_per_out[44]),
    .y_in(stage_3_per_out[45]),
    .x_out(stage_4_per_in[44]),
    .y_out(stage_4_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 68136911, 21713495, 7055647, 148662095, 256040960, 123185272, 170227406,
              193371292, 159404461, 183348420, 173702965, 186592442, 243304319, 236144340, 189591954,
              254509489, 66148505, 118518376, 108810259, 67012048, 104174682, 155168409, 3883583,
              25569479, 120936039, 13519489, 132703565, 71933862, 180525688, 139555205, 171721518}))
  stage_4_butterfly_23 (
    .x_in(stage_3_per_out[46]),
    .y_in(stage_3_per_out[47]),
    .x_out(stage_4_per_in[46]),
    .y_out(stage_4_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 68136911, 21713495, 7055647, 148662095, 256040960, 123185272, 170227406,
              193371292, 159404461, 183348420, 173702965, 186592442, 243304319, 236144340, 189591954,
              254509489, 66148505, 118518376, 108810259, 67012048, 104174682, 155168409, 3883583,
              25569479, 120936039, 13519489, 132703565, 71933862, 180525688, 139555205, 171721518}))
  stage_4_butterfly_24 (
    .x_in(stage_3_per_out[48]),
    .y_in(stage_3_per_out[49]),
    .x_out(stage_4_per_in[48]),
    .y_out(stage_4_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 68136911, 21713495, 7055647, 148662095, 256040960, 123185272, 170227406,
              193371292, 159404461, 183348420, 173702965, 186592442, 243304319, 236144340, 189591954,
              254509489, 66148505, 118518376, 108810259, 67012048, 104174682, 155168409, 3883583,
              25569479, 120936039, 13519489, 132703565, 71933862, 180525688, 139555205, 171721518}))
  stage_4_butterfly_25 (
    .x_in(stage_3_per_out[50]),
    .y_in(stage_3_per_out[51]),
    .x_out(stage_4_per_in[50]),
    .y_out(stage_4_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 68136911, 21713495, 7055647, 148662095, 256040960, 123185272, 170227406,
              193371292, 159404461, 183348420, 173702965, 186592442, 243304319, 236144340, 189591954,
              254509489, 66148505, 118518376, 108810259, 67012048, 104174682, 155168409, 3883583,
              25569479, 120936039, 13519489, 132703565, 71933862, 180525688, 139555205, 171721518}))
  stage_4_butterfly_26 (
    .x_in(stage_3_per_out[52]),
    .y_in(stage_3_per_out[53]),
    .x_out(stage_4_per_in[52]),
    .y_out(stage_4_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 68136911, 21713495, 7055647, 148662095, 256040960, 123185272, 170227406,
              193371292, 159404461, 183348420, 173702965, 186592442, 243304319, 236144340, 189591954,
              254509489, 66148505, 118518376, 108810259, 67012048, 104174682, 155168409, 3883583,
              25569479, 120936039, 13519489, 132703565, 71933862, 180525688, 139555205, 171721518}))
  stage_4_butterfly_27 (
    .x_in(stage_3_per_out[54]),
    .y_in(stage_3_per_out[55]),
    .x_out(stage_4_per_in[54]),
    .y_out(stage_4_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 68136911, 21713495, 7055647, 148662095, 256040960, 123185272, 170227406,
              193371292, 159404461, 183348420, 173702965, 186592442, 243304319, 236144340, 189591954,
              254509489, 66148505, 118518376, 108810259, 67012048, 104174682, 155168409, 3883583,
              25569479, 120936039, 13519489, 132703565, 71933862, 180525688, 139555205, 171721518}))
  stage_4_butterfly_28 (
    .x_in(stage_3_per_out[56]),
    .y_in(stage_3_per_out[57]),
    .x_out(stage_4_per_in[56]),
    .y_out(stage_4_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 68136911, 21713495, 7055647, 148662095, 256040960, 123185272, 170227406,
              193371292, 159404461, 183348420, 173702965, 186592442, 243304319, 236144340, 189591954,
              254509489, 66148505, 118518376, 108810259, 67012048, 104174682, 155168409, 3883583,
              25569479, 120936039, 13519489, 132703565, 71933862, 180525688, 139555205, 171721518}))
  stage_4_butterfly_29 (
    .x_in(stage_3_per_out[58]),
    .y_in(stage_3_per_out[59]),
    .x_out(stage_4_per_in[58]),
    .y_out(stage_4_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 68136911, 21713495, 7055647, 148662095, 256040960, 123185272, 170227406,
              193371292, 159404461, 183348420, 173702965, 186592442, 243304319, 236144340, 189591954,
              254509489, 66148505, 118518376, 108810259, 67012048, 104174682, 155168409, 3883583,
              25569479, 120936039, 13519489, 132703565, 71933862, 180525688, 139555205, 171721518}))
  stage_4_butterfly_30 (
    .x_in(stage_3_per_out[60]),
    .y_in(stage_3_per_out[61]),
    .x_out(stage_4_per_in[60]),
    .y_out(stage_4_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({261793746, 68136911, 21713495, 7055647, 148662095, 256040960, 123185272, 170227406,
              193371292, 159404461, 183348420, 173702965, 186592442, 243304319, 236144340, 189591954,
              254509489, 66148505, 118518376, 108810259, 67012048, 104174682, 155168409, 3883583,
              25569479, 120936039, 13519489, 132703565, 71933862, 180525688, 139555205, 171721518}))
  stage_4_butterfly_31 (
    .x_in(stage_3_per_out[62]),
    .y_in(stage_3_per_out[63]),
    .x_out(stage_4_per_in[62]),
    .y_out(stage_4_per_in[63]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({116401819, 71064168, 81956368, 135288005, 216143425, 265950570, 254450415, 14542514,
              250166212, 130557622, 234030247, 209086118, 10130658, 176471684, 231358848, 63350037,
              47751177, 229216409, 204666342, 33479018, 34119889, 2795054, 96142103, 41086336,
              211668928, 197074908, 252442032, 9720223, 143969713, 245828202, 98878775, 217644581}))
  stage_4_butterfly_32 (
    .x_in(stage_3_per_out[64]),
    .y_in(stage_3_per_out[65]),
    .x_out(stage_4_per_in[64]),
    .y_out(stage_4_per_in[65]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({116401819, 71064168, 81956368, 135288005, 216143425, 265950570, 254450415, 14542514,
              250166212, 130557622, 234030247, 209086118, 10130658, 176471684, 231358848, 63350037,
              47751177, 229216409, 204666342, 33479018, 34119889, 2795054, 96142103, 41086336,
              211668928, 197074908, 252442032, 9720223, 143969713, 245828202, 98878775, 217644581}))
  stage_4_butterfly_33 (
    .x_in(stage_3_per_out[66]),
    .y_in(stage_3_per_out[67]),
    .x_out(stage_4_per_in[66]),
    .y_out(stage_4_per_in[67]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({116401819, 71064168, 81956368, 135288005, 216143425, 265950570, 254450415, 14542514,
              250166212, 130557622, 234030247, 209086118, 10130658, 176471684, 231358848, 63350037,
              47751177, 229216409, 204666342, 33479018, 34119889, 2795054, 96142103, 41086336,
              211668928, 197074908, 252442032, 9720223, 143969713, 245828202, 98878775, 217644581}))
  stage_4_butterfly_34 (
    .x_in(stage_3_per_out[68]),
    .y_in(stage_3_per_out[69]),
    .x_out(stage_4_per_in[68]),
    .y_out(stage_4_per_in[69]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({116401819, 71064168, 81956368, 135288005, 216143425, 265950570, 254450415, 14542514,
              250166212, 130557622, 234030247, 209086118, 10130658, 176471684, 231358848, 63350037,
              47751177, 229216409, 204666342, 33479018, 34119889, 2795054, 96142103, 41086336,
              211668928, 197074908, 252442032, 9720223, 143969713, 245828202, 98878775, 217644581}))
  stage_4_butterfly_35 (
    .x_in(stage_3_per_out[70]),
    .y_in(stage_3_per_out[71]),
    .x_out(stage_4_per_in[70]),
    .y_out(stage_4_per_in[71]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({116401819, 71064168, 81956368, 135288005, 216143425, 265950570, 254450415, 14542514,
              250166212, 130557622, 234030247, 209086118, 10130658, 176471684, 231358848, 63350037,
              47751177, 229216409, 204666342, 33479018, 34119889, 2795054, 96142103, 41086336,
              211668928, 197074908, 252442032, 9720223, 143969713, 245828202, 98878775, 217644581}))
  stage_4_butterfly_36 (
    .x_in(stage_3_per_out[72]),
    .y_in(stage_3_per_out[73]),
    .x_out(stage_4_per_in[72]),
    .y_out(stage_4_per_in[73]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({116401819, 71064168, 81956368, 135288005, 216143425, 265950570, 254450415, 14542514,
              250166212, 130557622, 234030247, 209086118, 10130658, 176471684, 231358848, 63350037,
              47751177, 229216409, 204666342, 33479018, 34119889, 2795054, 96142103, 41086336,
              211668928, 197074908, 252442032, 9720223, 143969713, 245828202, 98878775, 217644581}))
  stage_4_butterfly_37 (
    .x_in(stage_3_per_out[74]),
    .y_in(stage_3_per_out[75]),
    .x_out(stage_4_per_in[74]),
    .y_out(stage_4_per_in[75]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({116401819, 71064168, 81956368, 135288005, 216143425, 265950570, 254450415, 14542514,
              250166212, 130557622, 234030247, 209086118, 10130658, 176471684, 231358848, 63350037,
              47751177, 229216409, 204666342, 33479018, 34119889, 2795054, 96142103, 41086336,
              211668928, 197074908, 252442032, 9720223, 143969713, 245828202, 98878775, 217644581}))
  stage_4_butterfly_38 (
    .x_in(stage_3_per_out[76]),
    .y_in(stage_3_per_out[77]),
    .x_out(stage_4_per_in[76]),
    .y_out(stage_4_per_in[77]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({116401819, 71064168, 81956368, 135288005, 216143425, 265950570, 254450415, 14542514,
              250166212, 130557622, 234030247, 209086118, 10130658, 176471684, 231358848, 63350037,
              47751177, 229216409, 204666342, 33479018, 34119889, 2795054, 96142103, 41086336,
              211668928, 197074908, 252442032, 9720223, 143969713, 245828202, 98878775, 217644581}))
  stage_4_butterfly_39 (
    .x_in(stage_3_per_out[78]),
    .y_in(stage_3_per_out[79]),
    .x_out(stage_4_per_in[78]),
    .y_out(stage_4_per_in[79]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({116401819, 71064168, 81956368, 135288005, 216143425, 265950570, 254450415, 14542514,
              250166212, 130557622, 234030247, 209086118, 10130658, 176471684, 231358848, 63350037,
              47751177, 229216409, 204666342, 33479018, 34119889, 2795054, 96142103, 41086336,
              211668928, 197074908, 252442032, 9720223, 143969713, 245828202, 98878775, 217644581}))
  stage_4_butterfly_40 (
    .x_in(stage_3_per_out[80]),
    .y_in(stage_3_per_out[81]),
    .x_out(stage_4_per_in[80]),
    .y_out(stage_4_per_in[81]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({116401819, 71064168, 81956368, 135288005, 216143425, 265950570, 254450415, 14542514,
              250166212, 130557622, 234030247, 209086118, 10130658, 176471684, 231358848, 63350037,
              47751177, 229216409, 204666342, 33479018, 34119889, 2795054, 96142103, 41086336,
              211668928, 197074908, 252442032, 9720223, 143969713, 245828202, 98878775, 217644581}))
  stage_4_butterfly_41 (
    .x_in(stage_3_per_out[82]),
    .y_in(stage_3_per_out[83]),
    .x_out(stage_4_per_in[82]),
    .y_out(stage_4_per_in[83]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({116401819, 71064168, 81956368, 135288005, 216143425, 265950570, 254450415, 14542514,
              250166212, 130557622, 234030247, 209086118, 10130658, 176471684, 231358848, 63350037,
              47751177, 229216409, 204666342, 33479018, 34119889, 2795054, 96142103, 41086336,
              211668928, 197074908, 252442032, 9720223, 143969713, 245828202, 98878775, 217644581}))
  stage_4_butterfly_42 (
    .x_in(stage_3_per_out[84]),
    .y_in(stage_3_per_out[85]),
    .x_out(stage_4_per_in[84]),
    .y_out(stage_4_per_in[85]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({116401819, 71064168, 81956368, 135288005, 216143425, 265950570, 254450415, 14542514,
              250166212, 130557622, 234030247, 209086118, 10130658, 176471684, 231358848, 63350037,
              47751177, 229216409, 204666342, 33479018, 34119889, 2795054, 96142103, 41086336,
              211668928, 197074908, 252442032, 9720223, 143969713, 245828202, 98878775, 217644581}))
  stage_4_butterfly_43 (
    .x_in(stage_3_per_out[86]),
    .y_in(stage_3_per_out[87]),
    .x_out(stage_4_per_in[86]),
    .y_out(stage_4_per_in[87]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({116401819, 71064168, 81956368, 135288005, 216143425, 265950570, 254450415, 14542514,
              250166212, 130557622, 234030247, 209086118, 10130658, 176471684, 231358848, 63350037,
              47751177, 229216409, 204666342, 33479018, 34119889, 2795054, 96142103, 41086336,
              211668928, 197074908, 252442032, 9720223, 143969713, 245828202, 98878775, 217644581}))
  stage_4_butterfly_44 (
    .x_in(stage_3_per_out[88]),
    .y_in(stage_3_per_out[89]),
    .x_out(stage_4_per_in[88]),
    .y_out(stage_4_per_in[89]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({116401819, 71064168, 81956368, 135288005, 216143425, 265950570, 254450415, 14542514,
              250166212, 130557622, 234030247, 209086118, 10130658, 176471684, 231358848, 63350037,
              47751177, 229216409, 204666342, 33479018, 34119889, 2795054, 96142103, 41086336,
              211668928, 197074908, 252442032, 9720223, 143969713, 245828202, 98878775, 217644581}))
  stage_4_butterfly_45 (
    .x_in(stage_3_per_out[90]),
    .y_in(stage_3_per_out[91]),
    .x_out(stage_4_per_in[90]),
    .y_out(stage_4_per_in[91]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({116401819, 71064168, 81956368, 135288005, 216143425, 265950570, 254450415, 14542514,
              250166212, 130557622, 234030247, 209086118, 10130658, 176471684, 231358848, 63350037,
              47751177, 229216409, 204666342, 33479018, 34119889, 2795054, 96142103, 41086336,
              211668928, 197074908, 252442032, 9720223, 143969713, 245828202, 98878775, 217644581}))
  stage_4_butterfly_46 (
    .x_in(stage_3_per_out[92]),
    .y_in(stage_3_per_out[93]),
    .x_out(stage_4_per_in[92]),
    .y_out(stage_4_per_in[93]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({116401819, 71064168, 81956368, 135288005, 216143425, 265950570, 254450415, 14542514,
              250166212, 130557622, 234030247, 209086118, 10130658, 176471684, 231358848, 63350037,
              47751177, 229216409, 204666342, 33479018, 34119889, 2795054, 96142103, 41086336,
              211668928, 197074908, 252442032, 9720223, 143969713, 245828202, 98878775, 217644581}))
  stage_4_butterfly_47 (
    .x_in(stage_3_per_out[94]),
    .y_in(stage_3_per_out[95]),
    .x_out(stage_4_per_in[94]),
    .y_out(stage_4_per_in[95]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({18729522, 166886297, 176917280, 238498066, 181639510, 240677074, 97765534, 40475021,
              167885779, 37051834, 41155851, 258612781, 139182289, 83853696, 230433664, 54284329,
              15417588, 108083129, 241682233, 223427563, 77337691, 161827885, 118841873, 134866823,
              123954975, 210298252, 162031725, 19493867, 230702770, 13250338, 9446767, 249970613}))
  stage_4_butterfly_48 (
    .x_in(stage_3_per_out[96]),
    .y_in(stage_3_per_out[97]),
    .x_out(stage_4_per_in[96]),
    .y_out(stage_4_per_in[97]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({18729522, 166886297, 176917280, 238498066, 181639510, 240677074, 97765534, 40475021,
              167885779, 37051834, 41155851, 258612781, 139182289, 83853696, 230433664, 54284329,
              15417588, 108083129, 241682233, 223427563, 77337691, 161827885, 118841873, 134866823,
              123954975, 210298252, 162031725, 19493867, 230702770, 13250338, 9446767, 249970613}))
  stage_4_butterfly_49 (
    .x_in(stage_3_per_out[98]),
    .y_in(stage_3_per_out[99]),
    .x_out(stage_4_per_in[98]),
    .y_out(stage_4_per_in[99]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({18729522, 166886297, 176917280, 238498066, 181639510, 240677074, 97765534, 40475021,
              167885779, 37051834, 41155851, 258612781, 139182289, 83853696, 230433664, 54284329,
              15417588, 108083129, 241682233, 223427563, 77337691, 161827885, 118841873, 134866823,
              123954975, 210298252, 162031725, 19493867, 230702770, 13250338, 9446767, 249970613}))
  stage_4_butterfly_50 (
    .x_in(stage_3_per_out[100]),
    .y_in(stage_3_per_out[101]),
    .x_out(stage_4_per_in[100]),
    .y_out(stage_4_per_in[101]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({18729522, 166886297, 176917280, 238498066, 181639510, 240677074, 97765534, 40475021,
              167885779, 37051834, 41155851, 258612781, 139182289, 83853696, 230433664, 54284329,
              15417588, 108083129, 241682233, 223427563, 77337691, 161827885, 118841873, 134866823,
              123954975, 210298252, 162031725, 19493867, 230702770, 13250338, 9446767, 249970613}))
  stage_4_butterfly_51 (
    .x_in(stage_3_per_out[102]),
    .y_in(stage_3_per_out[103]),
    .x_out(stage_4_per_in[102]),
    .y_out(stage_4_per_in[103]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({18729522, 166886297, 176917280, 238498066, 181639510, 240677074, 97765534, 40475021,
              167885779, 37051834, 41155851, 258612781, 139182289, 83853696, 230433664, 54284329,
              15417588, 108083129, 241682233, 223427563, 77337691, 161827885, 118841873, 134866823,
              123954975, 210298252, 162031725, 19493867, 230702770, 13250338, 9446767, 249970613}))
  stage_4_butterfly_52 (
    .x_in(stage_3_per_out[104]),
    .y_in(stage_3_per_out[105]),
    .x_out(stage_4_per_in[104]),
    .y_out(stage_4_per_in[105]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({18729522, 166886297, 176917280, 238498066, 181639510, 240677074, 97765534, 40475021,
              167885779, 37051834, 41155851, 258612781, 139182289, 83853696, 230433664, 54284329,
              15417588, 108083129, 241682233, 223427563, 77337691, 161827885, 118841873, 134866823,
              123954975, 210298252, 162031725, 19493867, 230702770, 13250338, 9446767, 249970613}))
  stage_4_butterfly_53 (
    .x_in(stage_3_per_out[106]),
    .y_in(stage_3_per_out[107]),
    .x_out(stage_4_per_in[106]),
    .y_out(stage_4_per_in[107]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({18729522, 166886297, 176917280, 238498066, 181639510, 240677074, 97765534, 40475021,
              167885779, 37051834, 41155851, 258612781, 139182289, 83853696, 230433664, 54284329,
              15417588, 108083129, 241682233, 223427563, 77337691, 161827885, 118841873, 134866823,
              123954975, 210298252, 162031725, 19493867, 230702770, 13250338, 9446767, 249970613}))
  stage_4_butterfly_54 (
    .x_in(stage_3_per_out[108]),
    .y_in(stage_3_per_out[109]),
    .x_out(stage_4_per_in[108]),
    .y_out(stage_4_per_in[109]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({18729522, 166886297, 176917280, 238498066, 181639510, 240677074, 97765534, 40475021,
              167885779, 37051834, 41155851, 258612781, 139182289, 83853696, 230433664, 54284329,
              15417588, 108083129, 241682233, 223427563, 77337691, 161827885, 118841873, 134866823,
              123954975, 210298252, 162031725, 19493867, 230702770, 13250338, 9446767, 249970613}))
  stage_4_butterfly_55 (
    .x_in(stage_3_per_out[110]),
    .y_in(stage_3_per_out[111]),
    .x_out(stage_4_per_in[110]),
    .y_out(stage_4_per_in[111]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({18729522, 166886297, 176917280, 238498066, 181639510, 240677074, 97765534, 40475021,
              167885779, 37051834, 41155851, 258612781, 139182289, 83853696, 230433664, 54284329,
              15417588, 108083129, 241682233, 223427563, 77337691, 161827885, 118841873, 134866823,
              123954975, 210298252, 162031725, 19493867, 230702770, 13250338, 9446767, 249970613}))
  stage_4_butterfly_56 (
    .x_in(stage_3_per_out[112]),
    .y_in(stage_3_per_out[113]),
    .x_out(stage_4_per_in[112]),
    .y_out(stage_4_per_in[113]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({18729522, 166886297, 176917280, 238498066, 181639510, 240677074, 97765534, 40475021,
              167885779, 37051834, 41155851, 258612781, 139182289, 83853696, 230433664, 54284329,
              15417588, 108083129, 241682233, 223427563, 77337691, 161827885, 118841873, 134866823,
              123954975, 210298252, 162031725, 19493867, 230702770, 13250338, 9446767, 249970613}))
  stage_4_butterfly_57 (
    .x_in(stage_3_per_out[114]),
    .y_in(stage_3_per_out[115]),
    .x_out(stage_4_per_in[114]),
    .y_out(stage_4_per_in[115]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({18729522, 166886297, 176917280, 238498066, 181639510, 240677074, 97765534, 40475021,
              167885779, 37051834, 41155851, 258612781, 139182289, 83853696, 230433664, 54284329,
              15417588, 108083129, 241682233, 223427563, 77337691, 161827885, 118841873, 134866823,
              123954975, 210298252, 162031725, 19493867, 230702770, 13250338, 9446767, 249970613}))
  stage_4_butterfly_58 (
    .x_in(stage_3_per_out[116]),
    .y_in(stage_3_per_out[117]),
    .x_out(stage_4_per_in[116]),
    .y_out(stage_4_per_in[117]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({18729522, 166886297, 176917280, 238498066, 181639510, 240677074, 97765534, 40475021,
              167885779, 37051834, 41155851, 258612781, 139182289, 83853696, 230433664, 54284329,
              15417588, 108083129, 241682233, 223427563, 77337691, 161827885, 118841873, 134866823,
              123954975, 210298252, 162031725, 19493867, 230702770, 13250338, 9446767, 249970613}))
  stage_4_butterfly_59 (
    .x_in(stage_3_per_out[118]),
    .y_in(stage_3_per_out[119]),
    .x_out(stage_4_per_in[118]),
    .y_out(stage_4_per_in[119]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({18729522, 166886297, 176917280, 238498066, 181639510, 240677074, 97765534, 40475021,
              167885779, 37051834, 41155851, 258612781, 139182289, 83853696, 230433664, 54284329,
              15417588, 108083129, 241682233, 223427563, 77337691, 161827885, 118841873, 134866823,
              123954975, 210298252, 162031725, 19493867, 230702770, 13250338, 9446767, 249970613}))
  stage_4_butterfly_60 (
    .x_in(stage_3_per_out[120]),
    .y_in(stage_3_per_out[121]),
    .x_out(stage_4_per_in[120]),
    .y_out(stage_4_per_in[121]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({18729522, 166886297, 176917280, 238498066, 181639510, 240677074, 97765534, 40475021,
              167885779, 37051834, 41155851, 258612781, 139182289, 83853696, 230433664, 54284329,
              15417588, 108083129, 241682233, 223427563, 77337691, 161827885, 118841873, 134866823,
              123954975, 210298252, 162031725, 19493867, 230702770, 13250338, 9446767, 249970613}))
  stage_4_butterfly_61 (
    .x_in(stage_3_per_out[122]),
    .y_in(stage_3_per_out[123]),
    .x_out(stage_4_per_in[122]),
    .y_out(stage_4_per_in[123]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({18729522, 166886297, 176917280, 238498066, 181639510, 240677074, 97765534, 40475021,
              167885779, 37051834, 41155851, 258612781, 139182289, 83853696, 230433664, 54284329,
              15417588, 108083129, 241682233, 223427563, 77337691, 161827885, 118841873, 134866823,
              123954975, 210298252, 162031725, 19493867, 230702770, 13250338, 9446767, 249970613}))
  stage_4_butterfly_62 (
    .x_in(stage_3_per_out[124]),
    .y_in(stage_3_per_out[125]),
    .x_out(stage_4_per_in[124]),
    .y_out(stage_4_per_in[125]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({18729522, 166886297, 176917280, 238498066, 181639510, 240677074, 97765534, 40475021,
              167885779, 37051834, 41155851, 258612781, 139182289, 83853696, 230433664, 54284329,
              15417588, 108083129, 241682233, 223427563, 77337691, 161827885, 118841873, 134866823,
              123954975, 210298252, 162031725, 19493867, 230702770, 13250338, 9446767, 249970613}))
  stage_4_butterfly_63 (
    .x_in(stage_3_per_out[126]),
    .y_in(stage_3_per_out[127]),
    .x_out(stage_4_per_in[126]),
    .y_out(stage_4_per_in[127]),
    .clk(clk),
    .rst(rst)
  );




  // TODO(Yang): stage 4 -> stage 5 permutation
  // FIXME: ignore butterfly units for now.
  stage_4_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_4_5_per (
    .inData_0(stage_4_per_in[0]),
    .inData_1(stage_4_per_in[1]),
    .inData_2(stage_4_per_in[2]),
    .inData_3(stage_4_per_in[3]),
    .inData_4(stage_4_per_in[4]),
    .inData_5(stage_4_per_in[5]),
    .inData_6(stage_4_per_in[6]),
    .inData_7(stage_4_per_in[7]),
    .inData_8(stage_4_per_in[8]),
    .inData_9(stage_4_per_in[9]),
    .inData_10(stage_4_per_in[10]),
    .inData_11(stage_4_per_in[11]),
    .inData_12(stage_4_per_in[12]),
    .inData_13(stage_4_per_in[13]),
    .inData_14(stage_4_per_in[14]),
    .inData_15(stage_4_per_in[15]),
    .inData_16(stage_4_per_in[16]),
    .inData_17(stage_4_per_in[17]),
    .inData_18(stage_4_per_in[18]),
    .inData_19(stage_4_per_in[19]),
    .inData_20(stage_4_per_in[20]),
    .inData_21(stage_4_per_in[21]),
    .inData_22(stage_4_per_in[22]),
    .inData_23(stage_4_per_in[23]),
    .inData_24(stage_4_per_in[24]),
    .inData_25(stage_4_per_in[25]),
    .inData_26(stage_4_per_in[26]),
    .inData_27(stage_4_per_in[27]),
    .inData_28(stage_4_per_in[28]),
    .inData_29(stage_4_per_in[29]),
    .inData_30(stage_4_per_in[30]),
    .inData_31(stage_4_per_in[31]),
    .inData_32(stage_4_per_in[32]),
    .inData_33(stage_4_per_in[33]),
    .inData_34(stage_4_per_in[34]),
    .inData_35(stage_4_per_in[35]),
    .inData_36(stage_4_per_in[36]),
    .inData_37(stage_4_per_in[37]),
    .inData_38(stage_4_per_in[38]),
    .inData_39(stage_4_per_in[39]),
    .inData_40(stage_4_per_in[40]),
    .inData_41(stage_4_per_in[41]),
    .inData_42(stage_4_per_in[42]),
    .inData_43(stage_4_per_in[43]),
    .inData_44(stage_4_per_in[44]),
    .inData_45(stage_4_per_in[45]),
    .inData_46(stage_4_per_in[46]),
    .inData_47(stage_4_per_in[47]),
    .inData_48(stage_4_per_in[48]),
    .inData_49(stage_4_per_in[49]),
    .inData_50(stage_4_per_in[50]),
    .inData_51(stage_4_per_in[51]),
    .inData_52(stage_4_per_in[52]),
    .inData_53(stage_4_per_in[53]),
    .inData_54(stage_4_per_in[54]),
    .inData_55(stage_4_per_in[55]),
    .inData_56(stage_4_per_in[56]),
    .inData_57(stage_4_per_in[57]),
    .inData_58(stage_4_per_in[58]),
    .inData_59(stage_4_per_in[59]),
    .inData_60(stage_4_per_in[60]),
    .inData_61(stage_4_per_in[61]),
    .inData_62(stage_4_per_in[62]),
    .inData_63(stage_4_per_in[63]),
    .inData_64(stage_4_per_in[64]),
    .inData_65(stage_4_per_in[65]),
    .inData_66(stage_4_per_in[66]),
    .inData_67(stage_4_per_in[67]),
    .inData_68(stage_4_per_in[68]),
    .inData_69(stage_4_per_in[69]),
    .inData_70(stage_4_per_in[70]),
    .inData_71(stage_4_per_in[71]),
    .inData_72(stage_4_per_in[72]),
    .inData_73(stage_4_per_in[73]),
    .inData_74(stage_4_per_in[74]),
    .inData_75(stage_4_per_in[75]),
    .inData_76(stage_4_per_in[76]),
    .inData_77(stage_4_per_in[77]),
    .inData_78(stage_4_per_in[78]),
    .inData_79(stage_4_per_in[79]),
    .inData_80(stage_4_per_in[80]),
    .inData_81(stage_4_per_in[81]),
    .inData_82(stage_4_per_in[82]),
    .inData_83(stage_4_per_in[83]),
    .inData_84(stage_4_per_in[84]),
    .inData_85(stage_4_per_in[85]),
    .inData_86(stage_4_per_in[86]),
    .inData_87(stage_4_per_in[87]),
    .inData_88(stage_4_per_in[88]),
    .inData_89(stage_4_per_in[89]),
    .inData_90(stage_4_per_in[90]),
    .inData_91(stage_4_per_in[91]),
    .inData_92(stage_4_per_in[92]),
    .inData_93(stage_4_per_in[93]),
    .inData_94(stage_4_per_in[94]),
    .inData_95(stage_4_per_in[95]),
    .inData_96(stage_4_per_in[96]),
    .inData_97(stage_4_per_in[97]),
    .inData_98(stage_4_per_in[98]),
    .inData_99(stage_4_per_in[99]),
    .inData_100(stage_4_per_in[100]),
    .inData_101(stage_4_per_in[101]),
    .inData_102(stage_4_per_in[102]),
    .inData_103(stage_4_per_in[103]),
    .inData_104(stage_4_per_in[104]),
    .inData_105(stage_4_per_in[105]),
    .inData_106(stage_4_per_in[106]),
    .inData_107(stage_4_per_in[107]),
    .inData_108(stage_4_per_in[108]),
    .inData_109(stage_4_per_in[109]),
    .inData_110(stage_4_per_in[110]),
    .inData_111(stage_4_per_in[111]),
    .inData_112(stage_4_per_in[112]),
    .inData_113(stage_4_per_in[113]),
    .inData_114(stage_4_per_in[114]),
    .inData_115(stage_4_per_in[115]),
    .inData_116(stage_4_per_in[116]),
    .inData_117(stage_4_per_in[117]),
    .inData_118(stage_4_per_in[118]),
    .inData_119(stage_4_per_in[119]),
    .inData_120(stage_4_per_in[120]),
    .inData_121(stage_4_per_in[121]),
    .inData_122(stage_4_per_in[122]),
    .inData_123(stage_4_per_in[123]),
    .inData_124(stage_4_per_in[124]),
    .inData_125(stage_4_per_in[125]),
    .inData_126(stage_4_per_in[126]),
    .inData_127(stage_4_per_in[127]),
    .outData_0(stage_4_per_out[0]),
    .outData_1(stage_4_per_out[1]),
    .outData_2(stage_4_per_out[2]),
    .outData_3(stage_4_per_out[3]),
    .outData_4(stage_4_per_out[4]),
    .outData_5(stage_4_per_out[5]),
    .outData_6(stage_4_per_out[6]),
    .outData_7(stage_4_per_out[7]),
    .outData_8(stage_4_per_out[8]),
    .outData_9(stage_4_per_out[9]),
    .outData_10(stage_4_per_out[10]),
    .outData_11(stage_4_per_out[11]),
    .outData_12(stage_4_per_out[12]),
    .outData_13(stage_4_per_out[13]),
    .outData_14(stage_4_per_out[14]),
    .outData_15(stage_4_per_out[15]),
    .outData_16(stage_4_per_out[16]),
    .outData_17(stage_4_per_out[17]),
    .outData_18(stage_4_per_out[18]),
    .outData_19(stage_4_per_out[19]),
    .outData_20(stage_4_per_out[20]),
    .outData_21(stage_4_per_out[21]),
    .outData_22(stage_4_per_out[22]),
    .outData_23(stage_4_per_out[23]),
    .outData_24(stage_4_per_out[24]),
    .outData_25(stage_4_per_out[25]),
    .outData_26(stage_4_per_out[26]),
    .outData_27(stage_4_per_out[27]),
    .outData_28(stage_4_per_out[28]),
    .outData_29(stage_4_per_out[29]),
    .outData_30(stage_4_per_out[30]),
    .outData_31(stage_4_per_out[31]),
    .outData_32(stage_4_per_out[32]),
    .outData_33(stage_4_per_out[33]),
    .outData_34(stage_4_per_out[34]),
    .outData_35(stage_4_per_out[35]),
    .outData_36(stage_4_per_out[36]),
    .outData_37(stage_4_per_out[37]),
    .outData_38(stage_4_per_out[38]),
    .outData_39(stage_4_per_out[39]),
    .outData_40(stage_4_per_out[40]),
    .outData_41(stage_4_per_out[41]),
    .outData_42(stage_4_per_out[42]),
    .outData_43(stage_4_per_out[43]),
    .outData_44(stage_4_per_out[44]),
    .outData_45(stage_4_per_out[45]),
    .outData_46(stage_4_per_out[46]),
    .outData_47(stage_4_per_out[47]),
    .outData_48(stage_4_per_out[48]),
    .outData_49(stage_4_per_out[49]),
    .outData_50(stage_4_per_out[50]),
    .outData_51(stage_4_per_out[51]),
    .outData_52(stage_4_per_out[52]),
    .outData_53(stage_4_per_out[53]),
    .outData_54(stage_4_per_out[54]),
    .outData_55(stage_4_per_out[55]),
    .outData_56(stage_4_per_out[56]),
    .outData_57(stage_4_per_out[57]),
    .outData_58(stage_4_per_out[58]),
    .outData_59(stage_4_per_out[59]),
    .outData_60(stage_4_per_out[60]),
    .outData_61(stage_4_per_out[61]),
    .outData_62(stage_4_per_out[62]),
    .outData_63(stage_4_per_out[63]),
    .outData_64(stage_4_per_out[64]),
    .outData_65(stage_4_per_out[65]),
    .outData_66(stage_4_per_out[66]),
    .outData_67(stage_4_per_out[67]),
    .outData_68(stage_4_per_out[68]),
    .outData_69(stage_4_per_out[69]),
    .outData_70(stage_4_per_out[70]),
    .outData_71(stage_4_per_out[71]),
    .outData_72(stage_4_per_out[72]),
    .outData_73(stage_4_per_out[73]),
    .outData_74(stage_4_per_out[74]),
    .outData_75(stage_4_per_out[75]),
    .outData_76(stage_4_per_out[76]),
    .outData_77(stage_4_per_out[77]),
    .outData_78(stage_4_per_out[78]),
    .outData_79(stage_4_per_out[79]),
    .outData_80(stage_4_per_out[80]),
    .outData_81(stage_4_per_out[81]),
    .outData_82(stage_4_per_out[82]),
    .outData_83(stage_4_per_out[83]),
    .outData_84(stage_4_per_out[84]),
    .outData_85(stage_4_per_out[85]),
    .outData_86(stage_4_per_out[86]),
    .outData_87(stage_4_per_out[87]),
    .outData_88(stage_4_per_out[88]),
    .outData_89(stage_4_per_out[89]),
    .outData_90(stage_4_per_out[90]),
    .outData_91(stage_4_per_out[91]),
    .outData_92(stage_4_per_out[92]),
    .outData_93(stage_4_per_out[93]),
    .outData_94(stage_4_per_out[94]),
    .outData_95(stage_4_per_out[95]),
    .outData_96(stage_4_per_out[96]),
    .outData_97(stage_4_per_out[97]),
    .outData_98(stage_4_per_out[98]),
    .outData_99(stage_4_per_out[99]),
    .outData_100(stage_4_per_out[100]),
    .outData_101(stage_4_per_out[101]),
    .outData_102(stage_4_per_out[102]),
    .outData_103(stage_4_per_out[103]),
    .outData_104(stage_4_per_out[104]),
    .outData_105(stage_4_per_out[105]),
    .outData_106(stage_4_per_out[106]),
    .outData_107(stage_4_per_out[107]),
    .outData_108(stage_4_per_out[108]),
    .outData_109(stage_4_per_out[109]),
    .outData_110(stage_4_per_out[110]),
    .outData_111(stage_4_per_out[111]),
    .outData_112(stage_4_per_out[112]),
    .outData_113(stage_4_per_out[113]),
    .outData_114(stage_4_per_out[114]),
    .outData_115(stage_4_per_out[115]),
    .outData_116(stage_4_per_out[116]),
    .outData_117(stage_4_per_out[117]),
    .outData_118(stage_4_per_out[118]),
    .outData_119(stage_4_per_out[119]),
    .outData_120(stage_4_per_out[120]),
    .outData_121(stage_4_per_out[121]),
    .outData_122(stage_4_per_out[122]),
    .outData_123(stage_4_per_out[123]),
    .outData_124(stage_4_per_out[124]),
    .outData_125(stage_4_per_out[125]),
    .outData_126(stage_4_per_out[126]),
    .outData_127(stage_4_per_out[127]),
    .in_start(in_start[4]),
    .out_start(out_start[4]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 5 32 butterfly units
  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_0 (
    .x_in(stage_4_per_out[0]),
    .y_in(stage_4_per_out[1]),
    .x_out(stage_5_per_in[0]),
    .y_out(stage_5_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_1 (
    .x_in(stage_4_per_out[2]),
    .y_in(stage_4_per_out[3]),
    .x_out(stage_5_per_in[2]),
    .y_out(stage_5_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_2 (
    .x_in(stage_4_per_out[4]),
    .y_in(stage_4_per_out[5]),
    .x_out(stage_5_per_in[4]),
    .y_out(stage_5_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_3 (
    .x_in(stage_4_per_out[6]),
    .y_in(stage_4_per_out[7]),
    .x_out(stage_5_per_in[6]),
    .y_out(stage_5_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_4 (
    .x_in(stage_4_per_out[8]),
    .y_in(stage_4_per_out[9]),
    .x_out(stage_5_per_in[8]),
    .y_out(stage_5_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_5 (
    .x_in(stage_4_per_out[10]),
    .y_in(stage_4_per_out[11]),
    .x_out(stage_5_per_in[10]),
    .y_out(stage_5_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_6 (
    .x_in(stage_4_per_out[12]),
    .y_in(stage_4_per_out[13]),
    .x_out(stage_5_per_in[12]),
    .y_out(stage_5_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_7 (
    .x_in(stage_4_per_out[14]),
    .y_in(stage_4_per_out[15]),
    .x_out(stage_5_per_in[14]),
    .y_out(stage_5_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_8 (
    .x_in(stage_4_per_out[16]),
    .y_in(stage_4_per_out[17]),
    .x_out(stage_5_per_in[16]),
    .y_out(stage_5_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_9 (
    .x_in(stage_4_per_out[18]),
    .y_in(stage_4_per_out[19]),
    .x_out(stage_5_per_in[18]),
    .y_out(stage_5_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_10 (
    .x_in(stage_4_per_out[20]),
    .y_in(stage_4_per_out[21]),
    .x_out(stage_5_per_in[20]),
    .y_out(stage_5_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_11 (
    .x_in(stage_4_per_out[22]),
    .y_in(stage_4_per_out[23]),
    .x_out(stage_5_per_in[22]),
    .y_out(stage_5_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_12 (
    .x_in(stage_4_per_out[24]),
    .y_in(stage_4_per_out[25]),
    .x_out(stage_5_per_in[24]),
    .y_out(stage_5_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_13 (
    .x_in(stage_4_per_out[26]),
    .y_in(stage_4_per_out[27]),
    .x_out(stage_5_per_in[26]),
    .y_out(stage_5_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_14 (
    .x_in(stage_4_per_out[28]),
    .y_in(stage_4_per_out[29]),
    .x_out(stage_5_per_in[28]),
    .y_out(stage_5_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_15 (
    .x_in(stage_4_per_out[30]),
    .y_in(stage_4_per_out[31]),
    .x_out(stage_5_per_in[30]),
    .y_out(stage_5_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_16 (
    .x_in(stage_4_per_out[32]),
    .y_in(stage_4_per_out[33]),
    .x_out(stage_5_per_in[32]),
    .y_out(stage_5_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_17 (
    .x_in(stage_4_per_out[34]),
    .y_in(stage_4_per_out[35]),
    .x_out(stage_5_per_in[34]),
    .y_out(stage_5_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_18 (
    .x_in(stage_4_per_out[36]),
    .y_in(stage_4_per_out[37]),
    .x_out(stage_5_per_in[36]),
    .y_out(stage_5_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_19 (
    .x_in(stage_4_per_out[38]),
    .y_in(stage_4_per_out[39]),
    .x_out(stage_5_per_in[38]),
    .y_out(stage_5_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_20 (
    .x_in(stage_4_per_out[40]),
    .y_in(stage_4_per_out[41]),
    .x_out(stage_5_per_in[40]),
    .y_out(stage_5_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_21 (
    .x_in(stage_4_per_out[42]),
    .y_in(stage_4_per_out[43]),
    .x_out(stage_5_per_in[42]),
    .y_out(stage_5_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_22 (
    .x_in(stage_4_per_out[44]),
    .y_in(stage_4_per_out[45]),
    .x_out(stage_5_per_in[44]),
    .y_out(stage_5_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_23 (
    .x_in(stage_4_per_out[46]),
    .y_in(stage_4_per_out[47]),
    .x_out(stage_5_per_in[46]),
    .y_out(stage_5_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_24 (
    .x_in(stage_4_per_out[48]),
    .y_in(stage_4_per_out[49]),
    .x_out(stage_5_per_in[48]),
    .y_out(stage_5_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_25 (
    .x_in(stage_4_per_out[50]),
    .y_in(stage_4_per_out[51]),
    .x_out(stage_5_per_in[50]),
    .y_out(stage_5_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_26 (
    .x_in(stage_4_per_out[52]),
    .y_in(stage_4_per_out[53]),
    .x_out(stage_5_per_in[52]),
    .y_out(stage_5_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_27 (
    .x_in(stage_4_per_out[54]),
    .y_in(stage_4_per_out[55]),
    .x_out(stage_5_per_in[54]),
    .y_out(stage_5_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_28 (
    .x_in(stage_4_per_out[56]),
    .y_in(stage_4_per_out[57]),
    .x_out(stage_5_per_in[56]),
    .y_out(stage_5_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_29 (
    .x_in(stage_4_per_out[58]),
    .y_in(stage_4_per_out[59]),
    .x_out(stage_5_per_in[58]),
    .y_out(stage_5_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_30 (
    .x_in(stage_4_per_out[60]),
    .y_in(stage_4_per_out[61]),
    .x_out(stage_5_per_in[60]),
    .y_out(stage_5_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 239095400, 169276669, 197386970, 159115155, 102065274, 157028693, 210568560,
              74680748, 155896930, 100099056, 136571165, 149429971, 175609590, 201062854, 191727270,
              227611463, 49823188, 202366126, 120670867, 256674305, 233560477, 92577793, 172642311,
              251290023, 202257393, 240684902, 263678998, 200054106, 140204941, 109553202, 262046585}))
  stage_5_butterfly_31 (
    .x_in(stage_4_per_out[62]),
    .y_in(stage_4_per_out[63]),
    .x_out(stage_5_per_in[62]),
    .y_out(stage_5_per_in[63]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_32 (
    .x_in(stage_4_per_out[64]),
    .y_in(stage_4_per_out[65]),
    .x_out(stage_5_per_in[64]),
    .y_out(stage_5_per_in[65]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_33 (
    .x_in(stage_4_per_out[66]),
    .y_in(stage_4_per_out[67]),
    .x_out(stage_5_per_in[66]),
    .y_out(stage_5_per_in[67]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_34 (
    .x_in(stage_4_per_out[68]),
    .y_in(stage_4_per_out[69]),
    .x_out(stage_5_per_in[68]),
    .y_out(stage_5_per_in[69]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_35 (
    .x_in(stage_4_per_out[70]),
    .y_in(stage_4_per_out[71]),
    .x_out(stage_5_per_in[70]),
    .y_out(stage_5_per_in[71]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_36 (
    .x_in(stage_4_per_out[72]),
    .y_in(stage_4_per_out[73]),
    .x_out(stage_5_per_in[72]),
    .y_out(stage_5_per_in[73]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_37 (
    .x_in(stage_4_per_out[74]),
    .y_in(stage_4_per_out[75]),
    .x_out(stage_5_per_in[74]),
    .y_out(stage_5_per_in[75]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_38 (
    .x_in(stage_4_per_out[76]),
    .y_in(stage_4_per_out[77]),
    .x_out(stage_5_per_in[76]),
    .y_out(stage_5_per_in[77]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_39 (
    .x_in(stage_4_per_out[78]),
    .y_in(stage_4_per_out[79]),
    .x_out(stage_5_per_in[78]),
    .y_out(stage_5_per_in[79]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_40 (
    .x_in(stage_4_per_out[80]),
    .y_in(stage_4_per_out[81]),
    .x_out(stage_5_per_in[80]),
    .y_out(stage_5_per_in[81]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_41 (
    .x_in(stage_4_per_out[82]),
    .y_in(stage_4_per_out[83]),
    .x_out(stage_5_per_in[82]),
    .y_out(stage_5_per_in[83]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_42 (
    .x_in(stage_4_per_out[84]),
    .y_in(stage_4_per_out[85]),
    .x_out(stage_5_per_in[84]),
    .y_out(stage_5_per_in[85]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_43 (
    .x_in(stage_4_per_out[86]),
    .y_in(stage_4_per_out[87]),
    .x_out(stage_5_per_in[86]),
    .y_out(stage_5_per_in[87]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_44 (
    .x_in(stage_4_per_out[88]),
    .y_in(stage_4_per_out[89]),
    .x_out(stage_5_per_in[88]),
    .y_out(stage_5_per_in[89]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_45 (
    .x_in(stage_4_per_out[90]),
    .y_in(stage_4_per_out[91]),
    .x_out(stage_5_per_in[90]),
    .y_out(stage_5_per_in[91]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_46 (
    .x_in(stage_4_per_out[92]),
    .y_in(stage_4_per_out[93]),
    .x_out(stage_5_per_in[92]),
    .y_out(stage_5_per_in[93]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_47 (
    .x_in(stage_4_per_out[94]),
    .y_in(stage_4_per_out[95]),
    .x_out(stage_5_per_in[94]),
    .y_out(stage_5_per_in[95]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_48 (
    .x_in(stage_4_per_out[96]),
    .y_in(stage_4_per_out[97]),
    .x_out(stage_5_per_in[96]),
    .y_out(stage_5_per_in[97]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_49 (
    .x_in(stage_4_per_out[98]),
    .y_in(stage_4_per_out[99]),
    .x_out(stage_5_per_in[98]),
    .y_out(stage_5_per_in[99]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_50 (
    .x_in(stage_4_per_out[100]),
    .y_in(stage_4_per_out[101]),
    .x_out(stage_5_per_in[100]),
    .y_out(stage_5_per_in[101]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_51 (
    .x_in(stage_4_per_out[102]),
    .y_in(stage_4_per_out[103]),
    .x_out(stage_5_per_in[102]),
    .y_out(stage_5_per_in[103]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_52 (
    .x_in(stage_4_per_out[104]),
    .y_in(stage_4_per_out[105]),
    .x_out(stage_5_per_in[104]),
    .y_out(stage_5_per_in[105]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_53 (
    .x_in(stage_4_per_out[106]),
    .y_in(stage_4_per_out[107]),
    .x_out(stage_5_per_in[106]),
    .y_out(stage_5_per_in[107]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_54 (
    .x_in(stage_4_per_out[108]),
    .y_in(stage_4_per_out[109]),
    .x_out(stage_5_per_in[108]),
    .y_out(stage_5_per_in[109]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_55 (
    .x_in(stage_4_per_out[110]),
    .y_in(stage_4_per_out[111]),
    .x_out(stage_5_per_in[110]),
    .y_out(stage_5_per_in[111]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_56 (
    .x_in(stage_4_per_out[112]),
    .y_in(stage_4_per_out[113]),
    .x_out(stage_5_per_in[112]),
    .y_out(stage_5_per_in[113]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_57 (
    .x_in(stage_4_per_out[114]),
    .y_in(stage_4_per_out[115]),
    .x_out(stage_5_per_in[114]),
    .y_out(stage_5_per_in[115]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_58 (
    .x_in(stage_4_per_out[116]),
    .y_in(stage_4_per_out[117]),
    .x_out(stage_5_per_in[116]),
    .y_out(stage_5_per_in[117]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_59 (
    .x_in(stage_4_per_out[118]),
    .y_in(stage_4_per_out[119]),
    .x_out(stage_5_per_in[118]),
    .y_out(stage_5_per_in[119]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_60 (
    .x_in(stage_4_per_out[120]),
    .y_in(stage_4_per_out[121]),
    .x_out(stage_5_per_in[120]),
    .y_out(stage_5_per_in[121]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_61 (
    .x_in(stage_4_per_out[122]),
    .y_in(stage_4_per_out[123]),
    .x_out(stage_5_per_in[122]),
    .y_out(stage_5_per_in[123]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_62 (
    .x_in(stage_4_per_out[124]),
    .y_in(stage_4_per_out[125]),
    .x_out(stage_5_per_in[124]),
    .y_out(stage_5_per_in[125]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({185598009, 39593842, 141548072, 119224607, 208403048, 111284191, 30748955, 91114882,
              162373432, 145384235, 71471012, 33165861, 206324144, 152865265, 138074788, 41084242,
              196909902, 78852289, 146694818, 86517113, 114407843, 78462606, 70582130, 215696667,
              193045667, 242795574, 47317233, 152412548, 76707105, 170752771, 179817683, 165226744}))
  stage_5_butterfly_63 (
    .x_in(stage_4_per_out[126]),
    .y_in(stage_4_per_out[127]),
    .x_out(stage_5_per_in[126]),
    .y_out(stage_5_per_in[127]),
    .clk(clk),
    .rst(rst)
  );



  // TODO(Yang): stage 5 -> stage 6 permutation
  // FIXME: ignore butterfly units for now.
  stage_5_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_5_6_per (
    .inData_0(stage_5_per_in[0]),
    .inData_1(stage_5_per_in[1]),
    .inData_2(stage_5_per_in[2]),
    .inData_3(stage_5_per_in[3]),
    .inData_4(stage_5_per_in[4]),
    .inData_5(stage_5_per_in[5]),
    .inData_6(stage_5_per_in[6]),
    .inData_7(stage_5_per_in[7]),
    .inData_8(stage_5_per_in[8]),
    .inData_9(stage_5_per_in[9]),
    .inData_10(stage_5_per_in[10]),
    .inData_11(stage_5_per_in[11]),
    .inData_12(stage_5_per_in[12]),
    .inData_13(stage_5_per_in[13]),
    .inData_14(stage_5_per_in[14]),
    .inData_15(stage_5_per_in[15]),
    .inData_16(stage_5_per_in[16]),
    .inData_17(stage_5_per_in[17]),
    .inData_18(stage_5_per_in[18]),
    .inData_19(stage_5_per_in[19]),
    .inData_20(stage_5_per_in[20]),
    .inData_21(stage_5_per_in[21]),
    .inData_22(stage_5_per_in[22]),
    .inData_23(stage_5_per_in[23]),
    .inData_24(stage_5_per_in[24]),
    .inData_25(stage_5_per_in[25]),
    .inData_26(stage_5_per_in[26]),
    .inData_27(stage_5_per_in[27]),
    .inData_28(stage_5_per_in[28]),
    .inData_29(stage_5_per_in[29]),
    .inData_30(stage_5_per_in[30]),
    .inData_31(stage_5_per_in[31]),
    .inData_32(stage_5_per_in[32]),
    .inData_33(stage_5_per_in[33]),
    .inData_34(stage_5_per_in[34]),
    .inData_35(stage_5_per_in[35]),
    .inData_36(stage_5_per_in[36]),
    .inData_37(stage_5_per_in[37]),
    .inData_38(stage_5_per_in[38]),
    .inData_39(stage_5_per_in[39]),
    .inData_40(stage_5_per_in[40]),
    .inData_41(stage_5_per_in[41]),
    .inData_42(stage_5_per_in[42]),
    .inData_43(stage_5_per_in[43]),
    .inData_44(stage_5_per_in[44]),
    .inData_45(stage_5_per_in[45]),
    .inData_46(stage_5_per_in[46]),
    .inData_47(stage_5_per_in[47]),
    .inData_48(stage_5_per_in[48]),
    .inData_49(stage_5_per_in[49]),
    .inData_50(stage_5_per_in[50]),
    .inData_51(stage_5_per_in[51]),
    .inData_52(stage_5_per_in[52]),
    .inData_53(stage_5_per_in[53]),
    .inData_54(stage_5_per_in[54]),
    .inData_55(stage_5_per_in[55]),
    .inData_56(stage_5_per_in[56]),
    .inData_57(stage_5_per_in[57]),
    .inData_58(stage_5_per_in[58]),
    .inData_59(stage_5_per_in[59]),
    .inData_60(stage_5_per_in[60]),
    .inData_61(stage_5_per_in[61]),
    .inData_62(stage_5_per_in[62]),
    .inData_63(stage_5_per_in[63]),
    .inData_64(stage_5_per_in[64]),
    .inData_65(stage_5_per_in[65]),
    .inData_66(stage_5_per_in[66]),
    .inData_67(stage_5_per_in[67]),
    .inData_68(stage_5_per_in[68]),
    .inData_69(stage_5_per_in[69]),
    .inData_70(stage_5_per_in[70]),
    .inData_71(stage_5_per_in[71]),
    .inData_72(stage_5_per_in[72]),
    .inData_73(stage_5_per_in[73]),
    .inData_74(stage_5_per_in[74]),
    .inData_75(stage_5_per_in[75]),
    .inData_76(stage_5_per_in[76]),
    .inData_77(stage_5_per_in[77]),
    .inData_78(stage_5_per_in[78]),
    .inData_79(stage_5_per_in[79]),
    .inData_80(stage_5_per_in[80]),
    .inData_81(stage_5_per_in[81]),
    .inData_82(stage_5_per_in[82]),
    .inData_83(stage_5_per_in[83]),
    .inData_84(stage_5_per_in[84]),
    .inData_85(stage_5_per_in[85]),
    .inData_86(stage_5_per_in[86]),
    .inData_87(stage_5_per_in[87]),
    .inData_88(stage_5_per_in[88]),
    .inData_89(stage_5_per_in[89]),
    .inData_90(stage_5_per_in[90]),
    .inData_91(stage_5_per_in[91]),
    .inData_92(stage_5_per_in[92]),
    .inData_93(stage_5_per_in[93]),
    .inData_94(stage_5_per_in[94]),
    .inData_95(stage_5_per_in[95]),
    .inData_96(stage_5_per_in[96]),
    .inData_97(stage_5_per_in[97]),
    .inData_98(stage_5_per_in[98]),
    .inData_99(stage_5_per_in[99]),
    .inData_100(stage_5_per_in[100]),
    .inData_101(stage_5_per_in[101]),
    .inData_102(stage_5_per_in[102]),
    .inData_103(stage_5_per_in[103]),
    .inData_104(stage_5_per_in[104]),
    .inData_105(stage_5_per_in[105]),
    .inData_106(stage_5_per_in[106]),
    .inData_107(stage_5_per_in[107]),
    .inData_108(stage_5_per_in[108]),
    .inData_109(stage_5_per_in[109]),
    .inData_110(stage_5_per_in[110]),
    .inData_111(stage_5_per_in[111]),
    .inData_112(stage_5_per_in[112]),
    .inData_113(stage_5_per_in[113]),
    .inData_114(stage_5_per_in[114]),
    .inData_115(stage_5_per_in[115]),
    .inData_116(stage_5_per_in[116]),
    .inData_117(stage_5_per_in[117]),
    .inData_118(stage_5_per_in[118]),
    .inData_119(stage_5_per_in[119]),
    .inData_120(stage_5_per_in[120]),
    .inData_121(stage_5_per_in[121]),
    .inData_122(stage_5_per_in[122]),
    .inData_123(stage_5_per_in[123]),
    .inData_124(stage_5_per_in[124]),
    .inData_125(stage_5_per_in[125]),
    .inData_126(stage_5_per_in[126]),
    .inData_127(stage_5_per_in[127]),
    .outData_0(stage_5_per_out[0]),
    .outData_1(stage_5_per_out[1]),
    .outData_2(stage_5_per_out[2]),
    .outData_3(stage_5_per_out[3]),
    .outData_4(stage_5_per_out[4]),
    .outData_5(stage_5_per_out[5]),
    .outData_6(stage_5_per_out[6]),
    .outData_7(stage_5_per_out[7]),
    .outData_8(stage_5_per_out[8]),
    .outData_9(stage_5_per_out[9]),
    .outData_10(stage_5_per_out[10]),
    .outData_11(stage_5_per_out[11]),
    .outData_12(stage_5_per_out[12]),
    .outData_13(stage_5_per_out[13]),
    .outData_14(stage_5_per_out[14]),
    .outData_15(stage_5_per_out[15]),
    .outData_16(stage_5_per_out[16]),
    .outData_17(stage_5_per_out[17]),
    .outData_18(stage_5_per_out[18]),
    .outData_19(stage_5_per_out[19]),
    .outData_20(stage_5_per_out[20]),
    .outData_21(stage_5_per_out[21]),
    .outData_22(stage_5_per_out[22]),
    .outData_23(stage_5_per_out[23]),
    .outData_24(stage_5_per_out[24]),
    .outData_25(stage_5_per_out[25]),
    .outData_26(stage_5_per_out[26]),
    .outData_27(stage_5_per_out[27]),
    .outData_28(stage_5_per_out[28]),
    .outData_29(stage_5_per_out[29]),
    .outData_30(stage_5_per_out[30]),
    .outData_31(stage_5_per_out[31]),
    .outData_32(stage_5_per_out[32]),
    .outData_33(stage_5_per_out[33]),
    .outData_34(stage_5_per_out[34]),
    .outData_35(stage_5_per_out[35]),
    .outData_36(stage_5_per_out[36]),
    .outData_37(stage_5_per_out[37]),
    .outData_38(stage_5_per_out[38]),
    .outData_39(stage_5_per_out[39]),
    .outData_40(stage_5_per_out[40]),
    .outData_41(stage_5_per_out[41]),
    .outData_42(stage_5_per_out[42]),
    .outData_43(stage_5_per_out[43]),
    .outData_44(stage_5_per_out[44]),
    .outData_45(stage_5_per_out[45]),
    .outData_46(stage_5_per_out[46]),
    .outData_47(stage_5_per_out[47]),
    .outData_48(stage_5_per_out[48]),
    .outData_49(stage_5_per_out[49]),
    .outData_50(stage_5_per_out[50]),
    .outData_51(stage_5_per_out[51]),
    .outData_52(stage_5_per_out[52]),
    .outData_53(stage_5_per_out[53]),
    .outData_54(stage_5_per_out[54]),
    .outData_55(stage_5_per_out[55]),
    .outData_56(stage_5_per_out[56]),
    .outData_57(stage_5_per_out[57]),
    .outData_58(stage_5_per_out[58]),
    .outData_59(stage_5_per_out[59]),
    .outData_60(stage_5_per_out[60]),
    .outData_61(stage_5_per_out[61]),
    .outData_62(stage_5_per_out[62]),
    .outData_63(stage_5_per_out[63]),
    .outData_64(stage_5_per_out[64]),
    .outData_65(stage_5_per_out[65]),
    .outData_66(stage_5_per_out[66]),
    .outData_67(stage_5_per_out[67]),
    .outData_68(stage_5_per_out[68]),
    .outData_69(stage_5_per_out[69]),
    .outData_70(stage_5_per_out[70]),
    .outData_71(stage_5_per_out[71]),
    .outData_72(stage_5_per_out[72]),
    .outData_73(stage_5_per_out[73]),
    .outData_74(stage_5_per_out[74]),
    .outData_75(stage_5_per_out[75]),
    .outData_76(stage_5_per_out[76]),
    .outData_77(stage_5_per_out[77]),
    .outData_78(stage_5_per_out[78]),
    .outData_79(stage_5_per_out[79]),
    .outData_80(stage_5_per_out[80]),
    .outData_81(stage_5_per_out[81]),
    .outData_82(stage_5_per_out[82]),
    .outData_83(stage_5_per_out[83]),
    .outData_84(stage_5_per_out[84]),
    .outData_85(stage_5_per_out[85]),
    .outData_86(stage_5_per_out[86]),
    .outData_87(stage_5_per_out[87]),
    .outData_88(stage_5_per_out[88]),
    .outData_89(stage_5_per_out[89]),
    .outData_90(stage_5_per_out[90]),
    .outData_91(stage_5_per_out[91]),
    .outData_92(stage_5_per_out[92]),
    .outData_93(stage_5_per_out[93]),
    .outData_94(stage_5_per_out[94]),
    .outData_95(stage_5_per_out[95]),
    .outData_96(stage_5_per_out[96]),
    .outData_97(stage_5_per_out[97]),
    .outData_98(stage_5_per_out[98]),
    .outData_99(stage_5_per_out[99]),
    .outData_100(stage_5_per_out[100]),
    .outData_101(stage_5_per_out[101]),
    .outData_102(stage_5_per_out[102]),
    .outData_103(stage_5_per_out[103]),
    .outData_104(stage_5_per_out[104]),
    .outData_105(stage_5_per_out[105]),
    .outData_106(stage_5_per_out[106]),
    .outData_107(stage_5_per_out[107]),
    .outData_108(stage_5_per_out[108]),
    .outData_109(stage_5_per_out[109]),
    .outData_110(stage_5_per_out[110]),
    .outData_111(stage_5_per_out[111]),
    .outData_112(stage_5_per_out[112]),
    .outData_113(stage_5_per_out[113]),
    .outData_114(stage_5_per_out[114]),
    .outData_115(stage_5_per_out[115]),
    .outData_116(stage_5_per_out[116]),
    .outData_117(stage_5_per_out[117]),
    .outData_118(stage_5_per_out[118]),
    .outData_119(stage_5_per_out[119]),
    .outData_120(stage_5_per_out[120]),
    .outData_121(stage_5_per_out[121]),
    .outData_122(stage_5_per_out[122]),
    .outData_123(stage_5_per_out[123]),
    .outData_124(stage_5_per_out[124]),
    .outData_125(stage_5_per_out[125]),
    .outData_126(stage_5_per_out[126]),
    .outData_127(stage_5_per_out[127]),
    .in_start(in_start[5]),
    .out_start(out_start[5]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 6 32 butterfly units
  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_0 (
    .x_in(stage_5_per_out[0]),
    .y_in(stage_5_per_out[1]),
    .x_out(stage_6_per_in[0]),
    .y_out(stage_6_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_1 (
    .x_in(stage_5_per_out[2]),
    .y_in(stage_5_per_out[3]),
    .x_out(stage_6_per_in[2]),
    .y_out(stage_6_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_2 (
    .x_in(stage_5_per_out[4]),
    .y_in(stage_5_per_out[5]),
    .x_out(stage_6_per_in[4]),
    .y_out(stage_6_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_3 (
    .x_in(stage_5_per_out[6]),
    .y_in(stage_5_per_out[7]),
    .x_out(stage_6_per_in[6]),
    .y_out(stage_6_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_4 (
    .x_in(stage_5_per_out[8]),
    .y_in(stage_5_per_out[9]),
    .x_out(stage_6_per_in[8]),
    .y_out(stage_6_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_5 (
    .x_in(stage_5_per_out[10]),
    .y_in(stage_5_per_out[11]),
    .x_out(stage_6_per_in[10]),
    .y_out(stage_6_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_6 (
    .x_in(stage_5_per_out[12]),
    .y_in(stage_5_per_out[13]),
    .x_out(stage_6_per_in[12]),
    .y_out(stage_6_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_7 (
    .x_in(stage_5_per_out[14]),
    .y_in(stage_5_per_out[15]),
    .x_out(stage_6_per_in[14]),
    .y_out(stage_6_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_8 (
    .x_in(stage_5_per_out[16]),
    .y_in(stage_5_per_out[17]),
    .x_out(stage_6_per_in[16]),
    .y_out(stage_6_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_9 (
    .x_in(stage_5_per_out[18]),
    .y_in(stage_5_per_out[19]),
    .x_out(stage_6_per_in[18]),
    .y_out(stage_6_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_10 (
    .x_in(stage_5_per_out[20]),
    .y_in(stage_5_per_out[21]),
    .x_out(stage_6_per_in[20]),
    .y_out(stage_6_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_11 (
    .x_in(stage_5_per_out[22]),
    .y_in(stage_5_per_out[23]),
    .x_out(stage_6_per_in[22]),
    .y_out(stage_6_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_12 (
    .x_in(stage_5_per_out[24]),
    .y_in(stage_5_per_out[25]),
    .x_out(stage_6_per_in[24]),
    .y_out(stage_6_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_13 (
    .x_in(stage_5_per_out[26]),
    .y_in(stage_5_per_out[27]),
    .x_out(stage_6_per_in[26]),
    .y_out(stage_6_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_14 (
    .x_in(stage_5_per_out[28]),
    .y_in(stage_5_per_out[29]),
    .x_out(stage_6_per_in[28]),
    .y_out(stage_6_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_15 (
    .x_in(stage_5_per_out[30]),
    .y_in(stage_5_per_out[31]),
    .x_out(stage_6_per_in[30]),
    .y_out(stage_6_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_16 (
    .x_in(stage_5_per_out[32]),
    .y_in(stage_5_per_out[33]),
    .x_out(stage_6_per_in[32]),
    .y_out(stage_6_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_17 (
    .x_in(stage_5_per_out[34]),
    .y_in(stage_5_per_out[35]),
    .x_out(stage_6_per_in[34]),
    .y_out(stage_6_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_18 (
    .x_in(stage_5_per_out[36]),
    .y_in(stage_5_per_out[37]),
    .x_out(stage_6_per_in[36]),
    .y_out(stage_6_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_19 (
    .x_in(stage_5_per_out[38]),
    .y_in(stage_5_per_out[39]),
    .x_out(stage_6_per_in[38]),
    .y_out(stage_6_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_20 (
    .x_in(stage_5_per_out[40]),
    .y_in(stage_5_per_out[41]),
    .x_out(stage_6_per_in[40]),
    .y_out(stage_6_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_21 (
    .x_in(stage_5_per_out[42]),
    .y_in(stage_5_per_out[43]),
    .x_out(stage_6_per_in[42]),
    .y_out(stage_6_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_22 (
    .x_in(stage_5_per_out[44]),
    .y_in(stage_5_per_out[45]),
    .x_out(stage_6_per_in[44]),
    .y_out(stage_6_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_23 (
    .x_in(stage_5_per_out[46]),
    .y_in(stage_5_per_out[47]),
    .x_out(stage_6_per_in[46]),
    .y_out(stage_6_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_24 (
    .x_in(stage_5_per_out[48]),
    .y_in(stage_5_per_out[49]),
    .x_out(stage_6_per_in[48]),
    .y_out(stage_6_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_25 (
    .x_in(stage_5_per_out[50]),
    .y_in(stage_5_per_out[51]),
    .x_out(stage_6_per_in[50]),
    .y_out(stage_6_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_26 (
    .x_in(stage_5_per_out[52]),
    .y_in(stage_5_per_out[53]),
    .x_out(stage_6_per_in[52]),
    .y_out(stage_6_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_27 (
    .x_in(stage_5_per_out[54]),
    .y_in(stage_5_per_out[55]),
    .x_out(stage_6_per_in[54]),
    .y_out(stage_6_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_28 (
    .x_in(stage_5_per_out[56]),
    .y_in(stage_5_per_out[57]),
    .x_out(stage_6_per_in[56]),
    .y_out(stage_6_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_29 (
    .x_in(stage_5_per_out[58]),
    .y_in(stage_5_per_out[59]),
    .x_out(stage_6_per_in[58]),
    .y_out(stage_6_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_30 (
    .x_in(stage_5_per_out[60]),
    .y_in(stage_5_per_out[61]),
    .x_out(stage_6_per_in[60]),
    .y_out(stage_6_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_31 (
    .x_in(stage_5_per_out[62]),
    .y_in(stage_5_per_out[63]),
    .x_out(stage_6_per_in[62]),
    .y_out(stage_6_per_in[63]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_32 (
    .x_in(stage_5_per_out[64]),
    .y_in(stage_5_per_out[65]),
    .x_out(stage_6_per_in[64]),
    .y_out(stage_6_per_in[65]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_33 (
    .x_in(stage_5_per_out[66]),
    .y_in(stage_5_per_out[67]),
    .x_out(stage_6_per_in[66]),
    .y_out(stage_6_per_in[67]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_34 (
    .x_in(stage_5_per_out[68]),
    .y_in(stage_5_per_out[69]),
    .x_out(stage_6_per_in[68]),
    .y_out(stage_6_per_in[69]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_35 (
    .x_in(stage_5_per_out[70]),
    .y_in(stage_5_per_out[71]),
    .x_out(stage_6_per_in[70]),
    .y_out(stage_6_per_in[71]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_36 (
    .x_in(stage_5_per_out[72]),
    .y_in(stage_5_per_out[73]),
    .x_out(stage_6_per_in[72]),
    .y_out(stage_6_per_in[73]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_37 (
    .x_in(stage_5_per_out[74]),
    .y_in(stage_5_per_out[75]),
    .x_out(stage_6_per_in[74]),
    .y_out(stage_6_per_in[75]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_38 (
    .x_in(stage_5_per_out[76]),
    .y_in(stage_5_per_out[77]),
    .x_out(stage_6_per_in[76]),
    .y_out(stage_6_per_in[77]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_39 (
    .x_in(stage_5_per_out[78]),
    .y_in(stage_5_per_out[79]),
    .x_out(stage_6_per_in[78]),
    .y_out(stage_6_per_in[79]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_40 (
    .x_in(stage_5_per_out[80]),
    .y_in(stage_5_per_out[81]),
    .x_out(stage_6_per_in[80]),
    .y_out(stage_6_per_in[81]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_41 (
    .x_in(stage_5_per_out[82]),
    .y_in(stage_5_per_out[83]),
    .x_out(stage_6_per_in[82]),
    .y_out(stage_6_per_in[83]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_42 (
    .x_in(stage_5_per_out[84]),
    .y_in(stage_5_per_out[85]),
    .x_out(stage_6_per_in[84]),
    .y_out(stage_6_per_in[85]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_43 (
    .x_in(stage_5_per_out[86]),
    .y_in(stage_5_per_out[87]),
    .x_out(stage_6_per_in[86]),
    .y_out(stage_6_per_in[87]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_44 (
    .x_in(stage_5_per_out[88]),
    .y_in(stage_5_per_out[89]),
    .x_out(stage_6_per_in[88]),
    .y_out(stage_6_per_in[89]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_45 (
    .x_in(stage_5_per_out[90]),
    .y_in(stage_5_per_out[91]),
    .x_out(stage_6_per_in[90]),
    .y_out(stage_6_per_in[91]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_46 (
    .x_in(stage_5_per_out[92]),
    .y_in(stage_5_per_out[93]),
    .x_out(stage_6_per_in[92]),
    .y_out(stage_6_per_in[93]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_47 (
    .x_in(stage_5_per_out[94]),
    .y_in(stage_5_per_out[95]),
    .x_out(stage_6_per_in[94]),
    .y_out(stage_6_per_in[95]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_48 (
    .x_in(stage_5_per_out[96]),
    .y_in(stage_5_per_out[97]),
    .x_out(stage_6_per_in[96]),
    .y_out(stage_6_per_in[97]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_49 (
    .x_in(stage_5_per_out[98]),
    .y_in(stage_5_per_out[99]),
    .x_out(stage_6_per_in[98]),
    .y_out(stage_6_per_in[99]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_50 (
    .x_in(stage_5_per_out[100]),
    .y_in(stage_5_per_out[101]),
    .x_out(stage_6_per_in[100]),
    .y_out(stage_6_per_in[101]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_51 (
    .x_in(stage_5_per_out[102]),
    .y_in(stage_5_per_out[103]),
    .x_out(stage_6_per_in[102]),
    .y_out(stage_6_per_in[103]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_52 (
    .x_in(stage_5_per_out[104]),
    .y_in(stage_5_per_out[105]),
    .x_out(stage_6_per_in[104]),
    .y_out(stage_6_per_in[105]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_53 (
    .x_in(stage_5_per_out[106]),
    .y_in(stage_5_per_out[107]),
    .x_out(stage_6_per_in[106]),
    .y_out(stage_6_per_in[107]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_54 (
    .x_in(stage_5_per_out[108]),
    .y_in(stage_5_per_out[109]),
    .x_out(stage_6_per_in[108]),
    .y_out(stage_6_per_in[109]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_55 (
    .x_in(stage_5_per_out[110]),
    .y_in(stage_5_per_out[111]),
    .x_out(stage_6_per_in[110]),
    .y_out(stage_6_per_in[111]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_56 (
    .x_in(stage_5_per_out[112]),
    .y_in(stage_5_per_out[113]),
    .x_out(stage_6_per_in[112]),
    .y_out(stage_6_per_in[113]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_57 (
    .x_in(stage_5_per_out[114]),
    .y_in(stage_5_per_out[115]),
    .x_out(stage_6_per_in[114]),
    .y_out(stage_6_per_in[115]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_58 (
    .x_in(stage_5_per_out[116]),
    .y_in(stage_5_per_out[117]),
    .x_out(stage_6_per_in[116]),
    .y_out(stage_6_per_in[117]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_59 (
    .x_in(stage_5_per_out[118]),
    .y_in(stage_5_per_out[119]),
    .x_out(stage_6_per_in[118]),
    .y_out(stage_6_per_in[119]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_60 (
    .x_in(stage_5_per_out[120]),
    .y_in(stage_5_per_out[121]),
    .x_out(stage_6_per_in[120]),
    .y_out(stage_6_per_in[121]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_61 (
    .x_in(stage_5_per_out[122]),
    .y_in(stage_5_per_out[123]),
    .x_out(stage_6_per_in[122]),
    .y_out(stage_6_per_in[123]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_62 (
    .x_in(stage_5_per_out[124]),
    .y_in(stage_5_per_out[125]),
    .x_out(stage_6_per_in[124]),
    .y_out(stage_6_per_in[125]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 102773617, 210831626, 84893967, 119480423, 102579498, 129001811, 72061017,
              72052889, 73825164, 18533839, 168579404, 47877183, 184798272, 5258704, 92744225,
              221840088, 216372172, 231414272, 94135184, 89995519, 220656190, 183300662, 160020761,
              249274747, 62061822, 76573097, 35289455, 234642902, 229105823, 256670830, 143639106}))
  stage_6_butterfly_63 (
    .x_in(stage_5_per_out[126]),
    .y_in(stage_5_per_out[127]),
    .x_out(stage_6_per_in[126]),
    .y_out(stage_6_per_in[127]),
    .clk(clk),
    .rst(rst)
  );





  // TODO(Yang): stage 6 -> stage 7 permutation
  // FIXME: ignore butterfly units for now.
  stage_6_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_6_7_per (
    .inData_0(stage_6_per_in[0]),
    .inData_1(stage_6_per_in[1]),
    .inData_2(stage_6_per_in[2]),
    .inData_3(stage_6_per_in[3]),
    .inData_4(stage_6_per_in[4]),
    .inData_5(stage_6_per_in[5]),
    .inData_6(stage_6_per_in[6]),
    .inData_7(stage_6_per_in[7]),
    .inData_8(stage_6_per_in[8]),
    .inData_9(stage_6_per_in[9]),
    .inData_10(stage_6_per_in[10]),
    .inData_11(stage_6_per_in[11]),
    .inData_12(stage_6_per_in[12]),
    .inData_13(stage_6_per_in[13]),
    .inData_14(stage_6_per_in[14]),
    .inData_15(stage_6_per_in[15]),
    .inData_16(stage_6_per_in[16]),
    .inData_17(stage_6_per_in[17]),
    .inData_18(stage_6_per_in[18]),
    .inData_19(stage_6_per_in[19]),
    .inData_20(stage_6_per_in[20]),
    .inData_21(stage_6_per_in[21]),
    .inData_22(stage_6_per_in[22]),
    .inData_23(stage_6_per_in[23]),
    .inData_24(stage_6_per_in[24]),
    .inData_25(stage_6_per_in[25]),
    .inData_26(stage_6_per_in[26]),
    .inData_27(stage_6_per_in[27]),
    .inData_28(stage_6_per_in[28]),
    .inData_29(stage_6_per_in[29]),
    .inData_30(stage_6_per_in[30]),
    .inData_31(stage_6_per_in[31]),
    .inData_32(stage_6_per_in[32]),
    .inData_33(stage_6_per_in[33]),
    .inData_34(stage_6_per_in[34]),
    .inData_35(stage_6_per_in[35]),
    .inData_36(stage_6_per_in[36]),
    .inData_37(stage_6_per_in[37]),
    .inData_38(stage_6_per_in[38]),
    .inData_39(stage_6_per_in[39]),
    .inData_40(stage_6_per_in[40]),
    .inData_41(stage_6_per_in[41]),
    .inData_42(stage_6_per_in[42]),
    .inData_43(stage_6_per_in[43]),
    .inData_44(stage_6_per_in[44]),
    .inData_45(stage_6_per_in[45]),
    .inData_46(stage_6_per_in[46]),
    .inData_47(stage_6_per_in[47]),
    .inData_48(stage_6_per_in[48]),
    .inData_49(stage_6_per_in[49]),
    .inData_50(stage_6_per_in[50]),
    .inData_51(stage_6_per_in[51]),
    .inData_52(stage_6_per_in[52]),
    .inData_53(stage_6_per_in[53]),
    .inData_54(stage_6_per_in[54]),
    .inData_55(stage_6_per_in[55]),
    .inData_56(stage_6_per_in[56]),
    .inData_57(stage_6_per_in[57]),
    .inData_58(stage_6_per_in[58]),
    .inData_59(stage_6_per_in[59]),
    .inData_60(stage_6_per_in[60]),
    .inData_61(stage_6_per_in[61]),
    .inData_62(stage_6_per_in[62]),
    .inData_63(stage_6_per_in[63]),
    .inData_64(stage_6_per_in[64]),
    .inData_65(stage_6_per_in[65]),
    .inData_66(stage_6_per_in[66]),
    .inData_67(stage_6_per_in[67]),
    .inData_68(stage_6_per_in[68]),
    .inData_69(stage_6_per_in[69]),
    .inData_70(stage_6_per_in[70]),
    .inData_71(stage_6_per_in[71]),
    .inData_72(stage_6_per_in[72]),
    .inData_73(stage_6_per_in[73]),
    .inData_74(stage_6_per_in[74]),
    .inData_75(stage_6_per_in[75]),
    .inData_76(stage_6_per_in[76]),
    .inData_77(stage_6_per_in[77]),
    .inData_78(stage_6_per_in[78]),
    .inData_79(stage_6_per_in[79]),
    .inData_80(stage_6_per_in[80]),
    .inData_81(stage_6_per_in[81]),
    .inData_82(stage_6_per_in[82]),
    .inData_83(stage_6_per_in[83]),
    .inData_84(stage_6_per_in[84]),
    .inData_85(stage_6_per_in[85]),
    .inData_86(stage_6_per_in[86]),
    .inData_87(stage_6_per_in[87]),
    .inData_88(stage_6_per_in[88]),
    .inData_89(stage_6_per_in[89]),
    .inData_90(stage_6_per_in[90]),
    .inData_91(stage_6_per_in[91]),
    .inData_92(stage_6_per_in[92]),
    .inData_93(stage_6_per_in[93]),
    .inData_94(stage_6_per_in[94]),
    .inData_95(stage_6_per_in[95]),
    .inData_96(stage_6_per_in[96]),
    .inData_97(stage_6_per_in[97]),
    .inData_98(stage_6_per_in[98]),
    .inData_99(stage_6_per_in[99]),
    .inData_100(stage_6_per_in[100]),
    .inData_101(stage_6_per_in[101]),
    .inData_102(stage_6_per_in[102]),
    .inData_103(stage_6_per_in[103]),
    .inData_104(stage_6_per_in[104]),
    .inData_105(stage_6_per_in[105]),
    .inData_106(stage_6_per_in[106]),
    .inData_107(stage_6_per_in[107]),
    .inData_108(stage_6_per_in[108]),
    .inData_109(stage_6_per_in[109]),
    .inData_110(stage_6_per_in[110]),
    .inData_111(stage_6_per_in[111]),
    .inData_112(stage_6_per_in[112]),
    .inData_113(stage_6_per_in[113]),
    .inData_114(stage_6_per_in[114]),
    .inData_115(stage_6_per_in[115]),
    .inData_116(stage_6_per_in[116]),
    .inData_117(stage_6_per_in[117]),
    .inData_118(stage_6_per_in[118]),
    .inData_119(stage_6_per_in[119]),
    .inData_120(stage_6_per_in[120]),
    .inData_121(stage_6_per_in[121]),
    .inData_122(stage_6_per_in[122]),
    .inData_123(stage_6_per_in[123]),
    .inData_124(stage_6_per_in[124]),
    .inData_125(stage_6_per_in[125]),
    .inData_126(stage_6_per_in[126]),
    .inData_127(stage_6_per_in[127]),
    .outData_0(stage_6_per_out[0]),
    .outData_1(stage_6_per_out[1]),
    .outData_2(stage_6_per_out[2]),
    .outData_3(stage_6_per_out[3]),
    .outData_4(stage_6_per_out[4]),
    .outData_5(stage_6_per_out[5]),
    .outData_6(stage_6_per_out[6]),
    .outData_7(stage_6_per_out[7]),
    .outData_8(stage_6_per_out[8]),
    .outData_9(stage_6_per_out[9]),
    .outData_10(stage_6_per_out[10]),
    .outData_11(stage_6_per_out[11]),
    .outData_12(stage_6_per_out[12]),
    .outData_13(stage_6_per_out[13]),
    .outData_14(stage_6_per_out[14]),
    .outData_15(stage_6_per_out[15]),
    .outData_16(stage_6_per_out[16]),
    .outData_17(stage_6_per_out[17]),
    .outData_18(stage_6_per_out[18]),
    .outData_19(stage_6_per_out[19]),
    .outData_20(stage_6_per_out[20]),
    .outData_21(stage_6_per_out[21]),
    .outData_22(stage_6_per_out[22]),
    .outData_23(stage_6_per_out[23]),
    .outData_24(stage_6_per_out[24]),
    .outData_25(stage_6_per_out[25]),
    .outData_26(stage_6_per_out[26]),
    .outData_27(stage_6_per_out[27]),
    .outData_28(stage_6_per_out[28]),
    .outData_29(stage_6_per_out[29]),
    .outData_30(stage_6_per_out[30]),
    .outData_31(stage_6_per_out[31]),
    .outData_32(stage_6_per_out[32]),
    .outData_33(stage_6_per_out[33]),
    .outData_34(stage_6_per_out[34]),
    .outData_35(stage_6_per_out[35]),
    .outData_36(stage_6_per_out[36]),
    .outData_37(stage_6_per_out[37]),
    .outData_38(stage_6_per_out[38]),
    .outData_39(stage_6_per_out[39]),
    .outData_40(stage_6_per_out[40]),
    .outData_41(stage_6_per_out[41]),
    .outData_42(stage_6_per_out[42]),
    .outData_43(stage_6_per_out[43]),
    .outData_44(stage_6_per_out[44]),
    .outData_45(stage_6_per_out[45]),
    .outData_46(stage_6_per_out[46]),
    .outData_47(stage_6_per_out[47]),
    .outData_48(stage_6_per_out[48]),
    .outData_49(stage_6_per_out[49]),
    .outData_50(stage_6_per_out[50]),
    .outData_51(stage_6_per_out[51]),
    .outData_52(stage_6_per_out[52]),
    .outData_53(stage_6_per_out[53]),
    .outData_54(stage_6_per_out[54]),
    .outData_55(stage_6_per_out[55]),
    .outData_56(stage_6_per_out[56]),
    .outData_57(stage_6_per_out[57]),
    .outData_58(stage_6_per_out[58]),
    .outData_59(stage_6_per_out[59]),
    .outData_60(stage_6_per_out[60]),
    .outData_61(stage_6_per_out[61]),
    .outData_62(stage_6_per_out[62]),
    .outData_63(stage_6_per_out[63]),
    .outData_64(stage_6_per_out[64]),
    .outData_65(stage_6_per_out[65]),
    .outData_66(stage_6_per_out[66]),
    .outData_67(stage_6_per_out[67]),
    .outData_68(stage_6_per_out[68]),
    .outData_69(stage_6_per_out[69]),
    .outData_70(stage_6_per_out[70]),
    .outData_71(stage_6_per_out[71]),
    .outData_72(stage_6_per_out[72]),
    .outData_73(stage_6_per_out[73]),
    .outData_74(stage_6_per_out[74]),
    .outData_75(stage_6_per_out[75]),
    .outData_76(stage_6_per_out[76]),
    .outData_77(stage_6_per_out[77]),
    .outData_78(stage_6_per_out[78]),
    .outData_79(stage_6_per_out[79]),
    .outData_80(stage_6_per_out[80]),
    .outData_81(stage_6_per_out[81]),
    .outData_82(stage_6_per_out[82]),
    .outData_83(stage_6_per_out[83]),
    .outData_84(stage_6_per_out[84]),
    .outData_85(stage_6_per_out[85]),
    .outData_86(stage_6_per_out[86]),
    .outData_87(stage_6_per_out[87]),
    .outData_88(stage_6_per_out[88]),
    .outData_89(stage_6_per_out[89]),
    .outData_90(stage_6_per_out[90]),
    .outData_91(stage_6_per_out[91]),
    .outData_92(stage_6_per_out[92]),
    .outData_93(stage_6_per_out[93]),
    .outData_94(stage_6_per_out[94]),
    .outData_95(stage_6_per_out[95]),
    .outData_96(stage_6_per_out[96]),
    .outData_97(stage_6_per_out[97]),
    .outData_98(stage_6_per_out[98]),
    .outData_99(stage_6_per_out[99]),
    .outData_100(stage_6_per_out[100]),
    .outData_101(stage_6_per_out[101]),
    .outData_102(stage_6_per_out[102]),
    .outData_103(stage_6_per_out[103]),
    .outData_104(stage_6_per_out[104]),
    .outData_105(stage_6_per_out[105]),
    .outData_106(stage_6_per_out[106]),
    .outData_107(stage_6_per_out[107]),
    .outData_108(stage_6_per_out[108]),
    .outData_109(stage_6_per_out[109]),
    .outData_110(stage_6_per_out[110]),
    .outData_111(stage_6_per_out[111]),
    .outData_112(stage_6_per_out[112]),
    .outData_113(stage_6_per_out[113]),
    .outData_114(stage_6_per_out[114]),
    .outData_115(stage_6_per_out[115]),
    .outData_116(stage_6_per_out[116]),
    .outData_117(stage_6_per_out[117]),
    .outData_118(stage_6_per_out[118]),
    .outData_119(stage_6_per_out[119]),
    .outData_120(stage_6_per_out[120]),
    .outData_121(stage_6_per_out[121]),
    .outData_122(stage_6_per_out[122]),
    .outData_123(stage_6_per_out[123]),
    .outData_124(stage_6_per_out[124]),
    .outData_125(stage_6_per_out[125]),
    .outData_126(stage_6_per_out[126]),
    .outData_127(stage_6_per_out[127]),
    .in_start(in_start[6]),
    .out_start(out_start[6]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 7 32 butterfly units
  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_0 (
    .x_in(stage_6_per_out[0]),
    .y_in(stage_6_per_out[1]),
    .x_out(stage_7_per_in[0]),
    .y_out(stage_7_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_1 (
    .x_in(stage_6_per_out[2]),
    .y_in(stage_6_per_out[3]),
    .x_out(stage_7_per_in[2]),
    .y_out(stage_7_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_2 (
    .x_in(stage_6_per_out[4]),
    .y_in(stage_6_per_out[5]),
    .x_out(stage_7_per_in[4]),
    .y_out(stage_7_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_3 (
    .x_in(stage_6_per_out[6]),
    .y_in(stage_6_per_out[7]),
    .x_out(stage_7_per_in[6]),
    .y_out(stage_7_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_4 (
    .x_in(stage_6_per_out[8]),
    .y_in(stage_6_per_out[9]),
    .x_out(stage_7_per_in[8]),
    .y_out(stage_7_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_5 (
    .x_in(stage_6_per_out[10]),
    .y_in(stage_6_per_out[11]),
    .x_out(stage_7_per_in[10]),
    .y_out(stage_7_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_6 (
    .x_in(stage_6_per_out[12]),
    .y_in(stage_6_per_out[13]),
    .x_out(stage_7_per_in[12]),
    .y_out(stage_7_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_7 (
    .x_in(stage_6_per_out[14]),
    .y_in(stage_6_per_out[15]),
    .x_out(stage_7_per_in[14]),
    .y_out(stage_7_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_8 (
    .x_in(stage_6_per_out[16]),
    .y_in(stage_6_per_out[17]),
    .x_out(stage_7_per_in[16]),
    .y_out(stage_7_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_9 (
    .x_in(stage_6_per_out[18]),
    .y_in(stage_6_per_out[19]),
    .x_out(stage_7_per_in[18]),
    .y_out(stage_7_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_10 (
    .x_in(stage_6_per_out[20]),
    .y_in(stage_6_per_out[21]),
    .x_out(stage_7_per_in[20]),
    .y_out(stage_7_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_11 (
    .x_in(stage_6_per_out[22]),
    .y_in(stage_6_per_out[23]),
    .x_out(stage_7_per_in[22]),
    .y_out(stage_7_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_12 (
    .x_in(stage_6_per_out[24]),
    .y_in(stage_6_per_out[25]),
    .x_out(stage_7_per_in[24]),
    .y_out(stage_7_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_13 (
    .x_in(stage_6_per_out[26]),
    .y_in(stage_6_per_out[27]),
    .x_out(stage_7_per_in[26]),
    .y_out(stage_7_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_14 (
    .x_in(stage_6_per_out[28]),
    .y_in(stage_6_per_out[29]),
    .x_out(stage_7_per_in[28]),
    .y_out(stage_7_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_15 (
    .x_in(stage_6_per_out[30]),
    .y_in(stage_6_per_out[31]),
    .x_out(stage_7_per_in[30]),
    .y_out(stage_7_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_16 (
    .x_in(stage_6_per_out[32]),
    .y_in(stage_6_per_out[33]),
    .x_out(stage_7_per_in[32]),
    .y_out(stage_7_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_17 (
    .x_in(stage_6_per_out[34]),
    .y_in(stage_6_per_out[35]),
    .x_out(stage_7_per_in[34]),
    .y_out(stage_7_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_18 (
    .x_in(stage_6_per_out[36]),
    .y_in(stage_6_per_out[37]),
    .x_out(stage_7_per_in[36]),
    .y_out(stage_7_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_19 (
    .x_in(stage_6_per_out[38]),
    .y_in(stage_6_per_out[39]),
    .x_out(stage_7_per_in[38]),
    .y_out(stage_7_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_20 (
    .x_in(stage_6_per_out[40]),
    .y_in(stage_6_per_out[41]),
    .x_out(stage_7_per_in[40]),
    .y_out(stage_7_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_21 (
    .x_in(stage_6_per_out[42]),
    .y_in(stage_6_per_out[43]),
    .x_out(stage_7_per_in[42]),
    .y_out(stage_7_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_22 (
    .x_in(stage_6_per_out[44]),
    .y_in(stage_6_per_out[45]),
    .x_out(stage_7_per_in[44]),
    .y_out(stage_7_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_23 (
    .x_in(stage_6_per_out[46]),
    .y_in(stage_6_per_out[47]),
    .x_out(stage_7_per_in[46]),
    .y_out(stage_7_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_24 (
    .x_in(stage_6_per_out[48]),
    .y_in(stage_6_per_out[49]),
    .x_out(stage_7_per_in[48]),
    .y_out(stage_7_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_25 (
    .x_in(stage_6_per_out[50]),
    .y_in(stage_6_per_out[51]),
    .x_out(stage_7_per_in[50]),
    .y_out(stage_7_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_26 (
    .x_in(stage_6_per_out[52]),
    .y_in(stage_6_per_out[53]),
    .x_out(stage_7_per_in[52]),
    .y_out(stage_7_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_27 (
    .x_in(stage_6_per_out[54]),
    .y_in(stage_6_per_out[55]),
    .x_out(stage_7_per_in[54]),
    .y_out(stage_7_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_28 (
    .x_in(stage_6_per_out[56]),
    .y_in(stage_6_per_out[57]),
    .x_out(stage_7_per_in[56]),
    .y_out(stage_7_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_29 (
    .x_in(stage_6_per_out[58]),
    .y_in(stage_6_per_out[59]),
    .x_out(stage_7_per_in[58]),
    .y_out(stage_7_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_30 (
    .x_in(stage_6_per_out[60]),
    .y_in(stage_6_per_out[61]),
    .x_out(stage_7_per_in[60]),
    .y_out(stage_7_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_31 (
    .x_in(stage_6_per_out[62]),
    .y_in(stage_6_per_out[63]),
    .x_out(stage_7_per_in[62]),
    .y_out(stage_7_per_in[63]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_32 (
    .x_in(stage_6_per_out[64]),
    .y_in(stage_6_per_out[65]),
    .x_out(stage_7_per_in[64]),
    .y_out(stage_7_per_in[65]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_33 (
    .x_in(stage_6_per_out[66]),
    .y_in(stage_6_per_out[67]),
    .x_out(stage_7_per_in[66]),
    .y_out(stage_7_per_in[67]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_34 (
    .x_in(stage_6_per_out[68]),
    .y_in(stage_6_per_out[69]),
    .x_out(stage_7_per_in[68]),
    .y_out(stage_7_per_in[69]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_35 (
    .x_in(stage_6_per_out[70]),
    .y_in(stage_6_per_out[71]),
    .x_out(stage_7_per_in[70]),
    .y_out(stage_7_per_in[71]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_36 (
    .x_in(stage_6_per_out[72]),
    .y_in(stage_6_per_out[73]),
    .x_out(stage_7_per_in[72]),
    .y_out(stage_7_per_in[73]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_37 (
    .x_in(stage_6_per_out[74]),
    .y_in(stage_6_per_out[75]),
    .x_out(stage_7_per_in[74]),
    .y_out(stage_7_per_in[75]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_38 (
    .x_in(stage_6_per_out[76]),
    .y_in(stage_6_per_out[77]),
    .x_out(stage_7_per_in[76]),
    .y_out(stage_7_per_in[77]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_39 (
    .x_in(stage_6_per_out[78]),
    .y_in(stage_6_per_out[79]),
    .x_out(stage_7_per_in[78]),
    .y_out(stage_7_per_in[79]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_40 (
    .x_in(stage_6_per_out[80]),
    .y_in(stage_6_per_out[81]),
    .x_out(stage_7_per_in[80]),
    .y_out(stage_7_per_in[81]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_41 (
    .x_in(stage_6_per_out[82]),
    .y_in(stage_6_per_out[83]),
    .x_out(stage_7_per_in[82]),
    .y_out(stage_7_per_in[83]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_42 (
    .x_in(stage_6_per_out[84]),
    .y_in(stage_6_per_out[85]),
    .x_out(stage_7_per_in[84]),
    .y_out(stage_7_per_in[85]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_43 (
    .x_in(stage_6_per_out[86]),
    .y_in(stage_6_per_out[87]),
    .x_out(stage_7_per_in[86]),
    .y_out(stage_7_per_in[87]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_44 (
    .x_in(stage_6_per_out[88]),
    .y_in(stage_6_per_out[89]),
    .x_out(stage_7_per_in[88]),
    .y_out(stage_7_per_in[89]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_45 (
    .x_in(stage_6_per_out[90]),
    .y_in(stage_6_per_out[91]),
    .x_out(stage_7_per_in[90]),
    .y_out(stage_7_per_in[91]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_46 (
    .x_in(stage_6_per_out[92]),
    .y_in(stage_6_per_out[93]),
    .x_out(stage_7_per_in[92]),
    .y_out(stage_7_per_in[93]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_47 (
    .x_in(stage_6_per_out[94]),
    .y_in(stage_6_per_out[95]),
    .x_out(stage_7_per_in[94]),
    .y_out(stage_7_per_in[95]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_48 (
    .x_in(stage_6_per_out[96]),
    .y_in(stage_6_per_out[97]),
    .x_out(stage_7_per_in[96]),
    .y_out(stage_7_per_in[97]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_49 (
    .x_in(stage_6_per_out[98]),
    .y_in(stage_6_per_out[99]),
    .x_out(stage_7_per_in[98]),
    .y_out(stage_7_per_in[99]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_50 (
    .x_in(stage_6_per_out[100]),
    .y_in(stage_6_per_out[101]),
    .x_out(stage_7_per_in[100]),
    .y_out(stage_7_per_in[101]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_51 (
    .x_in(stage_6_per_out[102]),
    .y_in(stage_6_per_out[103]),
    .x_out(stage_7_per_in[102]),
    .y_out(stage_7_per_in[103]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_52 (
    .x_in(stage_6_per_out[104]),
    .y_in(stage_6_per_out[105]),
    .x_out(stage_7_per_in[104]),
    .y_out(stage_7_per_in[105]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_53 (
    .x_in(stage_6_per_out[106]),
    .y_in(stage_6_per_out[107]),
    .x_out(stage_7_per_in[106]),
    .y_out(stage_7_per_in[107]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_54 (
    .x_in(stage_6_per_out[108]),
    .y_in(stage_6_per_out[109]),
    .x_out(stage_7_per_in[108]),
    .y_out(stage_7_per_in[109]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_55 (
    .x_in(stage_6_per_out[110]),
    .y_in(stage_6_per_out[111]),
    .x_out(stage_7_per_in[110]),
    .y_out(stage_7_per_in[111]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_56 (
    .x_in(stage_6_per_out[112]),
    .y_in(stage_6_per_out[113]),
    .x_out(stage_7_per_in[112]),
    .y_out(stage_7_per_in[113]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_57 (
    .x_in(stage_6_per_out[114]),
    .y_in(stage_6_per_out[115]),
    .x_out(stage_7_per_in[114]),
    .y_out(stage_7_per_in[115]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_58 (
    .x_in(stage_6_per_out[116]),
    .y_in(stage_6_per_out[117]),
    .x_out(stage_7_per_in[116]),
    .y_out(stage_7_per_in[117]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_59 (
    .x_in(stage_6_per_out[118]),
    .y_in(stage_6_per_out[119]),
    .x_out(stage_7_per_in[118]),
    .y_out(stage_7_per_in[119]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_60 (
    .x_in(stage_6_per_out[120]),
    .y_in(stage_6_per_out[121]),
    .x_out(stage_7_per_in[120]),
    .y_out(stage_7_per_in[121]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_61 (
    .x_in(stage_6_per_out[122]),
    .y_in(stage_6_per_out[123]),
    .x_out(stage_7_per_in[122]),
    .y_out(stage_7_per_in[123]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_62 (
    .x_in(stage_6_per_out[124]),
    .y_in(stage_6_per_out[125]),
    .x_out(stage_7_per_in[124]),
    .y_out(stage_7_per_in[125]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 33383981, 33383981, 125976015, 125976015, 69075086, 69075086,
              7802111, 7802111, 155624840, 155624840, 134587162, 134587162, 57620092, 57620092,
              133035932, 133035932, 225387856, 225387856, 163057267, 163057267, 73648196, 73648196,
              46265048, 46265048, 25800822, 25800822, 136955445, 136955445, 70516281, 70516281}))
  stage_7_butterfly_63 (
    .x_in(stage_6_per_out[126]),
    .y_in(stage_6_per_out[127]),
    .x_out(stage_7_per_in[126]),
    .y_out(stage_7_per_in[127]),
    .clk(clk),
    .rst(rst)
  );




  // TODO(Yang): stage 7 -> stage 8 permutation
  // FIXME: ignore butterfly units for now.
  stage_7_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_7_8_per (
    .inData_0(stage_7_per_in[0]),
    .inData_1(stage_7_per_in[1]),
    .inData_2(stage_7_per_in[2]),
    .inData_3(stage_7_per_in[3]),
    .inData_4(stage_7_per_in[4]),
    .inData_5(stage_7_per_in[5]),
    .inData_6(stage_7_per_in[6]),
    .inData_7(stage_7_per_in[7]),
    .inData_8(stage_7_per_in[8]),
    .inData_9(stage_7_per_in[9]),
    .inData_10(stage_7_per_in[10]),
    .inData_11(stage_7_per_in[11]),
    .inData_12(stage_7_per_in[12]),
    .inData_13(stage_7_per_in[13]),
    .inData_14(stage_7_per_in[14]),
    .inData_15(stage_7_per_in[15]),
    .inData_16(stage_7_per_in[16]),
    .inData_17(stage_7_per_in[17]),
    .inData_18(stage_7_per_in[18]),
    .inData_19(stage_7_per_in[19]),
    .inData_20(stage_7_per_in[20]),
    .inData_21(stage_7_per_in[21]),
    .inData_22(stage_7_per_in[22]),
    .inData_23(stage_7_per_in[23]),
    .inData_24(stage_7_per_in[24]),
    .inData_25(stage_7_per_in[25]),
    .inData_26(stage_7_per_in[26]),
    .inData_27(stage_7_per_in[27]),
    .inData_28(stage_7_per_in[28]),
    .inData_29(stage_7_per_in[29]),
    .inData_30(stage_7_per_in[30]),
    .inData_31(stage_7_per_in[31]),
    .inData_32(stage_7_per_in[32]),
    .inData_33(stage_7_per_in[33]),
    .inData_34(stage_7_per_in[34]),
    .inData_35(stage_7_per_in[35]),
    .inData_36(stage_7_per_in[36]),
    .inData_37(stage_7_per_in[37]),
    .inData_38(stage_7_per_in[38]),
    .inData_39(stage_7_per_in[39]),
    .inData_40(stage_7_per_in[40]),
    .inData_41(stage_7_per_in[41]),
    .inData_42(stage_7_per_in[42]),
    .inData_43(stage_7_per_in[43]),
    .inData_44(stage_7_per_in[44]),
    .inData_45(stage_7_per_in[45]),
    .inData_46(stage_7_per_in[46]),
    .inData_47(stage_7_per_in[47]),
    .inData_48(stage_7_per_in[48]),
    .inData_49(stage_7_per_in[49]),
    .inData_50(stage_7_per_in[50]),
    .inData_51(stage_7_per_in[51]),
    .inData_52(stage_7_per_in[52]),
    .inData_53(stage_7_per_in[53]),
    .inData_54(stage_7_per_in[54]),
    .inData_55(stage_7_per_in[55]),
    .inData_56(stage_7_per_in[56]),
    .inData_57(stage_7_per_in[57]),
    .inData_58(stage_7_per_in[58]),
    .inData_59(stage_7_per_in[59]),
    .inData_60(stage_7_per_in[60]),
    .inData_61(stage_7_per_in[61]),
    .inData_62(stage_7_per_in[62]),
    .inData_63(stage_7_per_in[63]),
    .inData_64(stage_7_per_in[64]),
    .inData_65(stage_7_per_in[65]),
    .inData_66(stage_7_per_in[66]),
    .inData_67(stage_7_per_in[67]),
    .inData_68(stage_7_per_in[68]),
    .inData_69(stage_7_per_in[69]),
    .inData_70(stage_7_per_in[70]),
    .inData_71(stage_7_per_in[71]),
    .inData_72(stage_7_per_in[72]),
    .inData_73(stage_7_per_in[73]),
    .inData_74(stage_7_per_in[74]),
    .inData_75(stage_7_per_in[75]),
    .inData_76(stage_7_per_in[76]),
    .inData_77(stage_7_per_in[77]),
    .inData_78(stage_7_per_in[78]),
    .inData_79(stage_7_per_in[79]),
    .inData_80(stage_7_per_in[80]),
    .inData_81(stage_7_per_in[81]),
    .inData_82(stage_7_per_in[82]),
    .inData_83(stage_7_per_in[83]),
    .inData_84(stage_7_per_in[84]),
    .inData_85(stage_7_per_in[85]),
    .inData_86(stage_7_per_in[86]),
    .inData_87(stage_7_per_in[87]),
    .inData_88(stage_7_per_in[88]),
    .inData_89(stage_7_per_in[89]),
    .inData_90(stage_7_per_in[90]),
    .inData_91(stage_7_per_in[91]),
    .inData_92(stage_7_per_in[92]),
    .inData_93(stage_7_per_in[93]),
    .inData_94(stage_7_per_in[94]),
    .inData_95(stage_7_per_in[95]),
    .inData_96(stage_7_per_in[96]),
    .inData_97(stage_7_per_in[97]),
    .inData_98(stage_7_per_in[98]),
    .inData_99(stage_7_per_in[99]),
    .inData_100(stage_7_per_in[100]),
    .inData_101(stage_7_per_in[101]),
    .inData_102(stage_7_per_in[102]),
    .inData_103(stage_7_per_in[103]),
    .inData_104(stage_7_per_in[104]),
    .inData_105(stage_7_per_in[105]),
    .inData_106(stage_7_per_in[106]),
    .inData_107(stage_7_per_in[107]),
    .inData_108(stage_7_per_in[108]),
    .inData_109(stage_7_per_in[109]),
    .inData_110(stage_7_per_in[110]),
    .inData_111(stage_7_per_in[111]),
    .inData_112(stage_7_per_in[112]),
    .inData_113(stage_7_per_in[113]),
    .inData_114(stage_7_per_in[114]),
    .inData_115(stage_7_per_in[115]),
    .inData_116(stage_7_per_in[116]),
    .inData_117(stage_7_per_in[117]),
    .inData_118(stage_7_per_in[118]),
    .inData_119(stage_7_per_in[119]),
    .inData_120(stage_7_per_in[120]),
    .inData_121(stage_7_per_in[121]),
    .inData_122(stage_7_per_in[122]),
    .inData_123(stage_7_per_in[123]),
    .inData_124(stage_7_per_in[124]),
    .inData_125(stage_7_per_in[125]),
    .inData_126(stage_7_per_in[126]),
    .inData_127(stage_7_per_in[127]),
    .outData_0(stage_7_per_out[0]),
    .outData_1(stage_7_per_out[1]),
    .outData_2(stage_7_per_out[2]),
    .outData_3(stage_7_per_out[3]),
    .outData_4(stage_7_per_out[4]),
    .outData_5(stage_7_per_out[5]),
    .outData_6(stage_7_per_out[6]),
    .outData_7(stage_7_per_out[7]),
    .outData_8(stage_7_per_out[8]),
    .outData_9(stage_7_per_out[9]),
    .outData_10(stage_7_per_out[10]),
    .outData_11(stage_7_per_out[11]),
    .outData_12(stage_7_per_out[12]),
    .outData_13(stage_7_per_out[13]),
    .outData_14(stage_7_per_out[14]),
    .outData_15(stage_7_per_out[15]),
    .outData_16(stage_7_per_out[16]),
    .outData_17(stage_7_per_out[17]),
    .outData_18(stage_7_per_out[18]),
    .outData_19(stage_7_per_out[19]),
    .outData_20(stage_7_per_out[20]),
    .outData_21(stage_7_per_out[21]),
    .outData_22(stage_7_per_out[22]),
    .outData_23(stage_7_per_out[23]),
    .outData_24(stage_7_per_out[24]),
    .outData_25(stage_7_per_out[25]),
    .outData_26(stage_7_per_out[26]),
    .outData_27(stage_7_per_out[27]),
    .outData_28(stage_7_per_out[28]),
    .outData_29(stage_7_per_out[29]),
    .outData_30(stage_7_per_out[30]),
    .outData_31(stage_7_per_out[31]),
    .outData_32(stage_7_per_out[32]),
    .outData_33(stage_7_per_out[33]),
    .outData_34(stage_7_per_out[34]),
    .outData_35(stage_7_per_out[35]),
    .outData_36(stage_7_per_out[36]),
    .outData_37(stage_7_per_out[37]),
    .outData_38(stage_7_per_out[38]),
    .outData_39(stage_7_per_out[39]),
    .outData_40(stage_7_per_out[40]),
    .outData_41(stage_7_per_out[41]),
    .outData_42(stage_7_per_out[42]),
    .outData_43(stage_7_per_out[43]),
    .outData_44(stage_7_per_out[44]),
    .outData_45(stage_7_per_out[45]),
    .outData_46(stage_7_per_out[46]),
    .outData_47(stage_7_per_out[47]),
    .outData_48(stage_7_per_out[48]),
    .outData_49(stage_7_per_out[49]),
    .outData_50(stage_7_per_out[50]),
    .outData_51(stage_7_per_out[51]),
    .outData_52(stage_7_per_out[52]),
    .outData_53(stage_7_per_out[53]),
    .outData_54(stage_7_per_out[54]),
    .outData_55(stage_7_per_out[55]),
    .outData_56(stage_7_per_out[56]),
    .outData_57(stage_7_per_out[57]),
    .outData_58(stage_7_per_out[58]),
    .outData_59(stage_7_per_out[59]),
    .outData_60(stage_7_per_out[60]),
    .outData_61(stage_7_per_out[61]),
    .outData_62(stage_7_per_out[62]),
    .outData_63(stage_7_per_out[63]),
    .outData_64(stage_7_per_out[64]),
    .outData_65(stage_7_per_out[65]),
    .outData_66(stage_7_per_out[66]),
    .outData_67(stage_7_per_out[67]),
    .outData_68(stage_7_per_out[68]),
    .outData_69(stage_7_per_out[69]),
    .outData_70(stage_7_per_out[70]),
    .outData_71(stage_7_per_out[71]),
    .outData_72(stage_7_per_out[72]),
    .outData_73(stage_7_per_out[73]),
    .outData_74(stage_7_per_out[74]),
    .outData_75(stage_7_per_out[75]),
    .outData_76(stage_7_per_out[76]),
    .outData_77(stage_7_per_out[77]),
    .outData_78(stage_7_per_out[78]),
    .outData_79(stage_7_per_out[79]),
    .outData_80(stage_7_per_out[80]),
    .outData_81(stage_7_per_out[81]),
    .outData_82(stage_7_per_out[82]),
    .outData_83(stage_7_per_out[83]),
    .outData_84(stage_7_per_out[84]),
    .outData_85(stage_7_per_out[85]),
    .outData_86(stage_7_per_out[86]),
    .outData_87(stage_7_per_out[87]),
    .outData_88(stage_7_per_out[88]),
    .outData_89(stage_7_per_out[89]),
    .outData_90(stage_7_per_out[90]),
    .outData_91(stage_7_per_out[91]),
    .outData_92(stage_7_per_out[92]),
    .outData_93(stage_7_per_out[93]),
    .outData_94(stage_7_per_out[94]),
    .outData_95(stage_7_per_out[95]),
    .outData_96(stage_7_per_out[96]),
    .outData_97(stage_7_per_out[97]),
    .outData_98(stage_7_per_out[98]),
    .outData_99(stage_7_per_out[99]),
    .outData_100(stage_7_per_out[100]),
    .outData_101(stage_7_per_out[101]),
    .outData_102(stage_7_per_out[102]),
    .outData_103(stage_7_per_out[103]),
    .outData_104(stage_7_per_out[104]),
    .outData_105(stage_7_per_out[105]),
    .outData_106(stage_7_per_out[106]),
    .outData_107(stage_7_per_out[107]),
    .outData_108(stage_7_per_out[108]),
    .outData_109(stage_7_per_out[109]),
    .outData_110(stage_7_per_out[110]),
    .outData_111(stage_7_per_out[111]),
    .outData_112(stage_7_per_out[112]),
    .outData_113(stage_7_per_out[113]),
    .outData_114(stage_7_per_out[114]),
    .outData_115(stage_7_per_out[115]),
    .outData_116(stage_7_per_out[116]),
    .outData_117(stage_7_per_out[117]),
    .outData_118(stage_7_per_out[118]),
    .outData_119(stage_7_per_out[119]),
    .outData_120(stage_7_per_out[120]),
    .outData_121(stage_7_per_out[121]),
    .outData_122(stage_7_per_out[122]),
    .outData_123(stage_7_per_out[123]),
    .outData_124(stage_7_per_out[124]),
    .outData_125(stage_7_per_out[125]),
    .outData_126(stage_7_per_out[126]),
    .outData_127(stage_7_per_out[127]),
    .in_start(in_start[7]),
    .out_start(out_start[7]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 8 32 butterfly units
  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_0 (
    .x_in(stage_7_per_out[0]),
    .y_in(stage_7_per_out[1]),
    .x_out(stage_8_per_in[0]),
    .y_out(stage_8_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_1 (
    .x_in(stage_7_per_out[2]),
    .y_in(stage_7_per_out[3]),
    .x_out(stage_8_per_in[2]),
    .y_out(stage_8_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_2 (
    .x_in(stage_7_per_out[4]),
    .y_in(stage_7_per_out[5]),
    .x_out(stage_8_per_in[4]),
    .y_out(stage_8_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_3 (
    .x_in(stage_7_per_out[6]),
    .y_in(stage_7_per_out[7]),
    .x_out(stage_8_per_in[6]),
    .y_out(stage_8_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_4 (
    .x_in(stage_7_per_out[8]),
    .y_in(stage_7_per_out[9]),
    .x_out(stage_8_per_in[8]),
    .y_out(stage_8_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_5 (
    .x_in(stage_7_per_out[10]),
    .y_in(stage_7_per_out[11]),
    .x_out(stage_8_per_in[10]),
    .y_out(stage_8_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_6 (
    .x_in(stage_7_per_out[12]),
    .y_in(stage_7_per_out[13]),
    .x_out(stage_8_per_in[12]),
    .y_out(stage_8_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_7 (
    .x_in(stage_7_per_out[14]),
    .y_in(stage_7_per_out[15]),
    .x_out(stage_8_per_in[14]),
    .y_out(stage_8_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_8 (
    .x_in(stage_7_per_out[16]),
    .y_in(stage_7_per_out[17]),
    .x_out(stage_8_per_in[16]),
    .y_out(stage_8_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_9 (
    .x_in(stage_7_per_out[18]),
    .y_in(stage_7_per_out[19]),
    .x_out(stage_8_per_in[18]),
    .y_out(stage_8_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_10 (
    .x_in(stage_7_per_out[20]),
    .y_in(stage_7_per_out[21]),
    .x_out(stage_8_per_in[20]),
    .y_out(stage_8_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_11 (
    .x_in(stage_7_per_out[22]),
    .y_in(stage_7_per_out[23]),
    .x_out(stage_8_per_in[22]),
    .y_out(stage_8_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_12 (
    .x_in(stage_7_per_out[24]),
    .y_in(stage_7_per_out[25]),
    .x_out(stage_8_per_in[24]),
    .y_out(stage_8_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_13 (
    .x_in(stage_7_per_out[26]),
    .y_in(stage_7_per_out[27]),
    .x_out(stage_8_per_in[26]),
    .y_out(stage_8_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_14 (
    .x_in(stage_7_per_out[28]),
    .y_in(stage_7_per_out[29]),
    .x_out(stage_8_per_in[28]),
    .y_out(stage_8_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_15 (
    .x_in(stage_7_per_out[30]),
    .y_in(stage_7_per_out[31]),
    .x_out(stage_8_per_in[30]),
    .y_out(stage_8_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_16 (
    .x_in(stage_7_per_out[32]),
    .y_in(stage_7_per_out[33]),
    .x_out(stage_8_per_in[32]),
    .y_out(stage_8_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_17 (
    .x_in(stage_7_per_out[34]),
    .y_in(stage_7_per_out[35]),
    .x_out(stage_8_per_in[34]),
    .y_out(stage_8_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_18 (
    .x_in(stage_7_per_out[36]),
    .y_in(stage_7_per_out[37]),
    .x_out(stage_8_per_in[36]),
    .y_out(stage_8_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_19 (
    .x_in(stage_7_per_out[38]),
    .y_in(stage_7_per_out[39]),
    .x_out(stage_8_per_in[38]),
    .y_out(stage_8_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_20 (
    .x_in(stage_7_per_out[40]),
    .y_in(stage_7_per_out[41]),
    .x_out(stage_8_per_in[40]),
    .y_out(stage_8_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_21 (
    .x_in(stage_7_per_out[42]),
    .y_in(stage_7_per_out[43]),
    .x_out(stage_8_per_in[42]),
    .y_out(stage_8_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_22 (
    .x_in(stage_7_per_out[44]),
    .y_in(stage_7_per_out[45]),
    .x_out(stage_8_per_in[44]),
    .y_out(stage_8_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_23 (
    .x_in(stage_7_per_out[46]),
    .y_in(stage_7_per_out[47]),
    .x_out(stage_8_per_in[46]),
    .y_out(stage_8_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_24 (
    .x_in(stage_7_per_out[48]),
    .y_in(stage_7_per_out[49]),
    .x_out(stage_8_per_in[48]),
    .y_out(stage_8_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_25 (
    .x_in(stage_7_per_out[50]),
    .y_in(stage_7_per_out[51]),
    .x_out(stage_8_per_in[50]),
    .y_out(stage_8_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_26 (
    .x_in(stage_7_per_out[52]),
    .y_in(stage_7_per_out[53]),
    .x_out(stage_8_per_in[52]),
    .y_out(stage_8_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_27 (
    .x_in(stage_7_per_out[54]),
    .y_in(stage_7_per_out[55]),
    .x_out(stage_8_per_in[54]),
    .y_out(stage_8_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_28 (
    .x_in(stage_7_per_out[56]),
    .y_in(stage_7_per_out[57]),
    .x_out(stage_8_per_in[56]),
    .y_out(stage_8_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_29 (
    .x_in(stage_7_per_out[58]),
    .y_in(stage_7_per_out[59]),
    .x_out(stage_8_per_in[58]),
    .y_out(stage_8_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_30 (
    .x_in(stage_7_per_out[60]),
    .y_in(stage_7_per_out[61]),
    .x_out(stage_8_per_in[60]),
    .y_out(stage_8_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_31 (
    .x_in(stage_7_per_out[62]),
    .y_in(stage_7_per_out[63]),
    .x_out(stage_8_per_in[62]),
    .y_out(stage_8_per_in[63]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_32 (
    .x_in(stage_7_per_out[64]),
    .y_in(stage_7_per_out[65]),
    .x_out(stage_8_per_in[64]),
    .y_out(stage_8_per_in[65]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_33 (
    .x_in(stage_7_per_out[66]),
    .y_in(stage_7_per_out[67]),
    .x_out(stage_8_per_in[66]),
    .y_out(stage_8_per_in[67]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_34 (
    .x_in(stage_7_per_out[68]),
    .y_in(stage_7_per_out[69]),
    .x_out(stage_8_per_in[68]),
    .y_out(stage_8_per_in[69]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_35 (
    .x_in(stage_7_per_out[70]),
    .y_in(stage_7_per_out[71]),
    .x_out(stage_8_per_in[70]),
    .y_out(stage_8_per_in[71]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_36 (
    .x_in(stage_7_per_out[72]),
    .y_in(stage_7_per_out[73]),
    .x_out(stage_8_per_in[72]),
    .y_out(stage_8_per_in[73]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_37 (
    .x_in(stage_7_per_out[74]),
    .y_in(stage_7_per_out[75]),
    .x_out(stage_8_per_in[74]),
    .y_out(stage_8_per_in[75]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_38 (
    .x_in(stage_7_per_out[76]),
    .y_in(stage_7_per_out[77]),
    .x_out(stage_8_per_in[76]),
    .y_out(stage_8_per_in[77]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_39 (
    .x_in(stage_7_per_out[78]),
    .y_in(stage_7_per_out[79]),
    .x_out(stage_8_per_in[78]),
    .y_out(stage_8_per_in[79]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_40 (
    .x_in(stage_7_per_out[80]),
    .y_in(stage_7_per_out[81]),
    .x_out(stage_8_per_in[80]),
    .y_out(stage_8_per_in[81]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_41 (
    .x_in(stage_7_per_out[82]),
    .y_in(stage_7_per_out[83]),
    .x_out(stage_8_per_in[82]),
    .y_out(stage_8_per_in[83]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_42 (
    .x_in(stage_7_per_out[84]),
    .y_in(stage_7_per_out[85]),
    .x_out(stage_8_per_in[84]),
    .y_out(stage_8_per_in[85]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_43 (
    .x_in(stage_7_per_out[86]),
    .y_in(stage_7_per_out[87]),
    .x_out(stage_8_per_in[86]),
    .y_out(stage_8_per_in[87]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_44 (
    .x_in(stage_7_per_out[88]),
    .y_in(stage_7_per_out[89]),
    .x_out(stage_8_per_in[88]),
    .y_out(stage_8_per_in[89]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_45 (
    .x_in(stage_7_per_out[90]),
    .y_in(stage_7_per_out[91]),
    .x_out(stage_8_per_in[90]),
    .y_out(stage_8_per_in[91]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_46 (
    .x_in(stage_7_per_out[92]),
    .y_in(stage_7_per_out[93]),
    .x_out(stage_8_per_in[92]),
    .y_out(stage_8_per_in[93]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_47 (
    .x_in(stage_7_per_out[94]),
    .y_in(stage_7_per_out[95]),
    .x_out(stage_8_per_in[94]),
    .y_out(stage_8_per_in[95]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_48 (
    .x_in(stage_7_per_out[96]),
    .y_in(stage_7_per_out[97]),
    .x_out(stage_8_per_in[96]),
    .y_out(stage_8_per_in[97]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_49 (
    .x_in(stage_7_per_out[98]),
    .y_in(stage_7_per_out[99]),
    .x_out(stage_8_per_in[98]),
    .y_out(stage_8_per_in[99]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_50 (
    .x_in(stage_7_per_out[100]),
    .y_in(stage_7_per_out[101]),
    .x_out(stage_8_per_in[100]),
    .y_out(stage_8_per_in[101]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_51 (
    .x_in(stage_7_per_out[102]),
    .y_in(stage_7_per_out[103]),
    .x_out(stage_8_per_in[102]),
    .y_out(stage_8_per_in[103]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_52 (
    .x_in(stage_7_per_out[104]),
    .y_in(stage_7_per_out[105]),
    .x_out(stage_8_per_in[104]),
    .y_out(stage_8_per_in[105]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_53 (
    .x_in(stage_7_per_out[106]),
    .y_in(stage_7_per_out[107]),
    .x_out(stage_8_per_in[106]),
    .y_out(stage_8_per_in[107]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_54 (
    .x_in(stage_7_per_out[108]),
    .y_in(stage_7_per_out[109]),
    .x_out(stage_8_per_in[108]),
    .y_out(stage_8_per_in[109]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_55 (
    .x_in(stage_7_per_out[110]),
    .y_in(stage_7_per_out[111]),
    .x_out(stage_8_per_in[110]),
    .y_out(stage_8_per_in[111]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_56 (
    .x_in(stage_7_per_out[112]),
    .y_in(stage_7_per_out[113]),
    .x_out(stage_8_per_in[112]),
    .y_out(stage_8_per_in[113]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_57 (
    .x_in(stage_7_per_out[114]),
    .y_in(stage_7_per_out[115]),
    .x_out(stage_8_per_in[114]),
    .y_out(stage_8_per_in[115]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_58 (
    .x_in(stage_7_per_out[116]),
    .y_in(stage_7_per_out[117]),
    .x_out(stage_8_per_in[116]),
    .y_out(stage_8_per_in[117]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_59 (
    .x_in(stage_7_per_out[118]),
    .y_in(stage_7_per_out[119]),
    .x_out(stage_8_per_in[118]),
    .y_out(stage_8_per_in[119]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_60 (
    .x_in(stage_7_per_out[120]),
    .y_in(stage_7_per_out[121]),
    .x_out(stage_8_per_in[120]),
    .y_out(stage_8_per_in[121]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_61 (
    .x_in(stage_7_per_out[122]),
    .y_in(stage_7_per_out[123]),
    .x_out(stage_8_per_in[122]),
    .y_out(stage_8_per_in[123]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_62 (
    .x_in(stage_7_per_out[124]),
    .y_in(stage_7_per_out[125]),
    .x_out(stage_8_per_in[124]),
    .y_out(stage_8_per_in[125]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_63 (
    .x_in(stage_7_per_out[126]),
    .y_in(stage_7_per_out[127]),
    .x_out(stage_8_per_in[126]),
    .y_out(stage_8_per_in[127]),
    .clk(clk),
    .rst(rst)
  );




  // TODO(Yang): stage 8 -> stage 9 permutation
  // FIXME: ignore butterfly units for now.
  stage_8_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_8_9_per (
    .inData_0(stage_8_per_in[0]),
    .inData_1(stage_8_per_in[1]),
    .inData_2(stage_8_per_in[2]),
    .inData_3(stage_8_per_in[3]),
    .inData_4(stage_8_per_in[4]),
    .inData_5(stage_8_per_in[5]),
    .inData_6(stage_8_per_in[6]),
    .inData_7(stage_8_per_in[7]),
    .inData_8(stage_8_per_in[8]),
    .inData_9(stage_8_per_in[9]),
    .inData_10(stage_8_per_in[10]),
    .inData_11(stage_8_per_in[11]),
    .inData_12(stage_8_per_in[12]),
    .inData_13(stage_8_per_in[13]),
    .inData_14(stage_8_per_in[14]),
    .inData_15(stage_8_per_in[15]),
    .inData_16(stage_8_per_in[16]),
    .inData_17(stage_8_per_in[17]),
    .inData_18(stage_8_per_in[18]),
    .inData_19(stage_8_per_in[19]),
    .inData_20(stage_8_per_in[20]),
    .inData_21(stage_8_per_in[21]),
    .inData_22(stage_8_per_in[22]),
    .inData_23(stage_8_per_in[23]),
    .inData_24(stage_8_per_in[24]),
    .inData_25(stage_8_per_in[25]),
    .inData_26(stage_8_per_in[26]),
    .inData_27(stage_8_per_in[27]),
    .inData_28(stage_8_per_in[28]),
    .inData_29(stage_8_per_in[29]),
    .inData_30(stage_8_per_in[30]),
    .inData_31(stage_8_per_in[31]),
    .inData_32(stage_8_per_in[32]),
    .inData_33(stage_8_per_in[33]),
    .inData_34(stage_8_per_in[34]),
    .inData_35(stage_8_per_in[35]),
    .inData_36(stage_8_per_in[36]),
    .inData_37(stage_8_per_in[37]),
    .inData_38(stage_8_per_in[38]),
    .inData_39(stage_8_per_in[39]),
    .inData_40(stage_8_per_in[40]),
    .inData_41(stage_8_per_in[41]),
    .inData_42(stage_8_per_in[42]),
    .inData_43(stage_8_per_in[43]),
    .inData_44(stage_8_per_in[44]),
    .inData_45(stage_8_per_in[45]),
    .inData_46(stage_8_per_in[46]),
    .inData_47(stage_8_per_in[47]),
    .inData_48(stage_8_per_in[48]),
    .inData_49(stage_8_per_in[49]),
    .inData_50(stage_8_per_in[50]),
    .inData_51(stage_8_per_in[51]),
    .inData_52(stage_8_per_in[52]),
    .inData_53(stage_8_per_in[53]),
    .inData_54(stage_8_per_in[54]),
    .inData_55(stage_8_per_in[55]),
    .inData_56(stage_8_per_in[56]),
    .inData_57(stage_8_per_in[57]),
    .inData_58(stage_8_per_in[58]),
    .inData_59(stage_8_per_in[59]),
    .inData_60(stage_8_per_in[60]),
    .inData_61(stage_8_per_in[61]),
    .inData_62(stage_8_per_in[62]),
    .inData_63(stage_8_per_in[63]),
    .inData_64(stage_8_per_in[64]),
    .inData_65(stage_8_per_in[65]),
    .inData_66(stage_8_per_in[66]),
    .inData_67(stage_8_per_in[67]),
    .inData_68(stage_8_per_in[68]),
    .inData_69(stage_8_per_in[69]),
    .inData_70(stage_8_per_in[70]),
    .inData_71(stage_8_per_in[71]),
    .inData_72(stage_8_per_in[72]),
    .inData_73(stage_8_per_in[73]),
    .inData_74(stage_8_per_in[74]),
    .inData_75(stage_8_per_in[75]),
    .inData_76(stage_8_per_in[76]),
    .inData_77(stage_8_per_in[77]),
    .inData_78(stage_8_per_in[78]),
    .inData_79(stage_8_per_in[79]),
    .inData_80(stage_8_per_in[80]),
    .inData_81(stage_8_per_in[81]),
    .inData_82(stage_8_per_in[82]),
    .inData_83(stage_8_per_in[83]),
    .inData_84(stage_8_per_in[84]),
    .inData_85(stage_8_per_in[85]),
    .inData_86(stage_8_per_in[86]),
    .inData_87(stage_8_per_in[87]),
    .inData_88(stage_8_per_in[88]),
    .inData_89(stage_8_per_in[89]),
    .inData_90(stage_8_per_in[90]),
    .inData_91(stage_8_per_in[91]),
    .inData_92(stage_8_per_in[92]),
    .inData_93(stage_8_per_in[93]),
    .inData_94(stage_8_per_in[94]),
    .inData_95(stage_8_per_in[95]),
    .inData_96(stage_8_per_in[96]),
    .inData_97(stage_8_per_in[97]),
    .inData_98(stage_8_per_in[98]),
    .inData_99(stage_8_per_in[99]),
    .inData_100(stage_8_per_in[100]),
    .inData_101(stage_8_per_in[101]),
    .inData_102(stage_8_per_in[102]),
    .inData_103(stage_8_per_in[103]),
    .inData_104(stage_8_per_in[104]),
    .inData_105(stage_8_per_in[105]),
    .inData_106(stage_8_per_in[106]),
    .inData_107(stage_8_per_in[107]),
    .inData_108(stage_8_per_in[108]),
    .inData_109(stage_8_per_in[109]),
    .inData_110(stage_8_per_in[110]),
    .inData_111(stage_8_per_in[111]),
    .inData_112(stage_8_per_in[112]),
    .inData_113(stage_8_per_in[113]),
    .inData_114(stage_8_per_in[114]),
    .inData_115(stage_8_per_in[115]),
    .inData_116(stage_8_per_in[116]),
    .inData_117(stage_8_per_in[117]),
    .inData_118(stage_8_per_in[118]),
    .inData_119(stage_8_per_in[119]),
    .inData_120(stage_8_per_in[120]),
    .inData_121(stage_8_per_in[121]),
    .inData_122(stage_8_per_in[122]),
    .inData_123(stage_8_per_in[123]),
    .inData_124(stage_8_per_in[124]),
    .inData_125(stage_8_per_in[125]),
    .inData_126(stage_8_per_in[126]),
    .inData_127(stage_8_per_in[127]),
    .outData_0(stage_8_per_out[0]),
    .outData_1(stage_8_per_out[1]),
    .outData_2(stage_8_per_out[2]),
    .outData_3(stage_8_per_out[3]),
    .outData_4(stage_8_per_out[4]),
    .outData_5(stage_8_per_out[5]),
    .outData_6(stage_8_per_out[6]),
    .outData_7(stage_8_per_out[7]),
    .outData_8(stage_8_per_out[8]),
    .outData_9(stage_8_per_out[9]),
    .outData_10(stage_8_per_out[10]),
    .outData_11(stage_8_per_out[11]),
    .outData_12(stage_8_per_out[12]),
    .outData_13(stage_8_per_out[13]),
    .outData_14(stage_8_per_out[14]),
    .outData_15(stage_8_per_out[15]),
    .outData_16(stage_8_per_out[16]),
    .outData_17(stage_8_per_out[17]),
    .outData_18(stage_8_per_out[18]),
    .outData_19(stage_8_per_out[19]),
    .outData_20(stage_8_per_out[20]),
    .outData_21(stage_8_per_out[21]),
    .outData_22(stage_8_per_out[22]),
    .outData_23(stage_8_per_out[23]),
    .outData_24(stage_8_per_out[24]),
    .outData_25(stage_8_per_out[25]),
    .outData_26(stage_8_per_out[26]),
    .outData_27(stage_8_per_out[27]),
    .outData_28(stage_8_per_out[28]),
    .outData_29(stage_8_per_out[29]),
    .outData_30(stage_8_per_out[30]),
    .outData_31(stage_8_per_out[31]),
    .outData_32(stage_8_per_out[32]),
    .outData_33(stage_8_per_out[33]),
    .outData_34(stage_8_per_out[34]),
    .outData_35(stage_8_per_out[35]),
    .outData_36(stage_8_per_out[36]),
    .outData_37(stage_8_per_out[37]),
    .outData_38(stage_8_per_out[38]),
    .outData_39(stage_8_per_out[39]),
    .outData_40(stage_8_per_out[40]),
    .outData_41(stage_8_per_out[41]),
    .outData_42(stage_8_per_out[42]),
    .outData_43(stage_8_per_out[43]),
    .outData_44(stage_8_per_out[44]),
    .outData_45(stage_8_per_out[45]),
    .outData_46(stage_8_per_out[46]),
    .outData_47(stage_8_per_out[47]),
    .outData_48(stage_8_per_out[48]),
    .outData_49(stage_8_per_out[49]),
    .outData_50(stage_8_per_out[50]),
    .outData_51(stage_8_per_out[51]),
    .outData_52(stage_8_per_out[52]),
    .outData_53(stage_8_per_out[53]),
    .outData_54(stage_8_per_out[54]),
    .outData_55(stage_8_per_out[55]),
    .outData_56(stage_8_per_out[56]),
    .outData_57(stage_8_per_out[57]),
    .outData_58(stage_8_per_out[58]),
    .outData_59(stage_8_per_out[59]),
    .outData_60(stage_8_per_out[60]),
    .outData_61(stage_8_per_out[61]),
    .outData_62(stage_8_per_out[62]),
    .outData_63(stage_8_per_out[63]),
    .outData_64(stage_8_per_out[64]),
    .outData_65(stage_8_per_out[65]),
    .outData_66(stage_8_per_out[66]),
    .outData_67(stage_8_per_out[67]),
    .outData_68(stage_8_per_out[68]),
    .outData_69(stage_8_per_out[69]),
    .outData_70(stage_8_per_out[70]),
    .outData_71(stage_8_per_out[71]),
    .outData_72(stage_8_per_out[72]),
    .outData_73(stage_8_per_out[73]),
    .outData_74(stage_8_per_out[74]),
    .outData_75(stage_8_per_out[75]),
    .outData_76(stage_8_per_out[76]),
    .outData_77(stage_8_per_out[77]),
    .outData_78(stage_8_per_out[78]),
    .outData_79(stage_8_per_out[79]),
    .outData_80(stage_8_per_out[80]),
    .outData_81(stage_8_per_out[81]),
    .outData_82(stage_8_per_out[82]),
    .outData_83(stage_8_per_out[83]),
    .outData_84(stage_8_per_out[84]),
    .outData_85(stage_8_per_out[85]),
    .outData_86(stage_8_per_out[86]),
    .outData_87(stage_8_per_out[87]),
    .outData_88(stage_8_per_out[88]),
    .outData_89(stage_8_per_out[89]),
    .outData_90(stage_8_per_out[90]),
    .outData_91(stage_8_per_out[91]),
    .outData_92(stage_8_per_out[92]),
    .outData_93(stage_8_per_out[93]),
    .outData_94(stage_8_per_out[94]),
    .outData_95(stage_8_per_out[95]),
    .outData_96(stage_8_per_out[96]),
    .outData_97(stage_8_per_out[97]),
    .outData_98(stage_8_per_out[98]),
    .outData_99(stage_8_per_out[99]),
    .outData_100(stage_8_per_out[100]),
    .outData_101(stage_8_per_out[101]),
    .outData_102(stage_8_per_out[102]),
    .outData_103(stage_8_per_out[103]),
    .outData_104(stage_8_per_out[104]),
    .outData_105(stage_8_per_out[105]),
    .outData_106(stage_8_per_out[106]),
    .outData_107(stage_8_per_out[107]),
    .outData_108(stage_8_per_out[108]),
    .outData_109(stage_8_per_out[109]),
    .outData_110(stage_8_per_out[110]),
    .outData_111(stage_8_per_out[111]),
    .outData_112(stage_8_per_out[112]),
    .outData_113(stage_8_per_out[113]),
    .outData_114(stage_8_per_out[114]),
    .outData_115(stage_8_per_out[115]),
    .outData_116(stage_8_per_out[116]),
    .outData_117(stage_8_per_out[117]),
    .outData_118(stage_8_per_out[118]),
    .outData_119(stage_8_per_out[119]),
    .outData_120(stage_8_per_out[120]),
    .outData_121(stage_8_per_out[121]),
    .outData_122(stage_8_per_out[122]),
    .outData_123(stage_8_per_out[123]),
    .outData_124(stage_8_per_out[124]),
    .outData_125(stage_8_per_out[125]),
    .outData_126(stage_8_per_out[126]),
    .outData_127(stage_8_per_out[127]),
    .in_start(in_start[8]),
    .out_start(out_start[8]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 9 32 butterfly units
  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_0 (
    .x_in(stage_8_per_out[0]),
    .y_in(stage_8_per_out[1]),
    .x_out(stage_9_per_in[0]),
    .y_out(stage_9_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_1 (
    .x_in(stage_8_per_out[2]),
    .y_in(stage_8_per_out[3]),
    .x_out(stage_9_per_in[2]),
    .y_out(stage_9_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_2 (
    .x_in(stage_8_per_out[4]),
    .y_in(stage_8_per_out[5]),
    .x_out(stage_9_per_in[4]),
    .y_out(stage_9_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_3 (
    .x_in(stage_8_per_out[6]),
    .y_in(stage_8_per_out[7]),
    .x_out(stage_9_per_in[6]),
    .y_out(stage_9_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_4 (
    .x_in(stage_8_per_out[8]),
    .y_in(stage_8_per_out[9]),
    .x_out(stage_9_per_in[8]),
    .y_out(stage_9_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_5 (
    .x_in(stage_8_per_out[10]),
    .y_in(stage_8_per_out[11]),
    .x_out(stage_9_per_in[10]),
    .y_out(stage_9_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_6 (
    .x_in(stage_8_per_out[12]),
    .y_in(stage_8_per_out[13]),
    .x_out(stage_9_per_in[12]),
    .y_out(stage_9_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_7 (
    .x_in(stage_8_per_out[14]),
    .y_in(stage_8_per_out[15]),
    .x_out(stage_9_per_in[14]),
    .y_out(stage_9_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_8 (
    .x_in(stage_8_per_out[16]),
    .y_in(stage_8_per_out[17]),
    .x_out(stage_9_per_in[16]),
    .y_out(stage_9_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_9 (
    .x_in(stage_8_per_out[18]),
    .y_in(stage_8_per_out[19]),
    .x_out(stage_9_per_in[18]),
    .y_out(stage_9_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_10 (
    .x_in(stage_8_per_out[20]),
    .y_in(stage_8_per_out[21]),
    .x_out(stage_9_per_in[20]),
    .y_out(stage_9_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_11 (
    .x_in(stage_8_per_out[22]),
    .y_in(stage_8_per_out[23]),
    .x_out(stage_9_per_in[22]),
    .y_out(stage_9_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_12 (
    .x_in(stage_8_per_out[24]),
    .y_in(stage_8_per_out[25]),
    .x_out(stage_9_per_in[24]),
    .y_out(stage_9_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_13 (
    .x_in(stage_8_per_out[26]),
    .y_in(stage_8_per_out[27]),
    .x_out(stage_9_per_in[26]),
    .y_out(stage_9_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_14 (
    .x_in(stage_8_per_out[28]),
    .y_in(stage_8_per_out[29]),
    .x_out(stage_9_per_in[28]),
    .y_out(stage_9_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_15 (
    .x_in(stage_8_per_out[30]),
    .y_in(stage_8_per_out[31]),
    .x_out(stage_9_per_in[30]),
    .y_out(stage_9_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_16 (
    .x_in(stage_8_per_out[32]),
    .y_in(stage_8_per_out[33]),
    .x_out(stage_9_per_in[32]),
    .y_out(stage_9_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_17 (
    .x_in(stage_8_per_out[34]),
    .y_in(stage_8_per_out[35]),
    .x_out(stage_9_per_in[34]),
    .y_out(stage_9_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_18 (
    .x_in(stage_8_per_out[36]),
    .y_in(stage_8_per_out[37]),
    .x_out(stage_9_per_in[36]),
    .y_out(stage_9_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_19 (
    .x_in(stage_8_per_out[38]),
    .y_in(stage_8_per_out[39]),
    .x_out(stage_9_per_in[38]),
    .y_out(stage_9_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_20 (
    .x_in(stage_8_per_out[40]),
    .y_in(stage_8_per_out[41]),
    .x_out(stage_9_per_in[40]),
    .y_out(stage_9_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_21 (
    .x_in(stage_8_per_out[42]),
    .y_in(stage_8_per_out[43]),
    .x_out(stage_9_per_in[42]),
    .y_out(stage_9_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_22 (
    .x_in(stage_8_per_out[44]),
    .y_in(stage_8_per_out[45]),
    .x_out(stage_9_per_in[44]),
    .y_out(stage_9_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_23 (
    .x_in(stage_8_per_out[46]),
    .y_in(stage_8_per_out[47]),
    .x_out(stage_9_per_in[46]),
    .y_out(stage_9_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_24 (
    .x_in(stage_8_per_out[48]),
    .y_in(stage_8_per_out[49]),
    .x_out(stage_9_per_in[48]),
    .y_out(stage_9_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_25 (
    .x_in(stage_8_per_out[50]),
    .y_in(stage_8_per_out[51]),
    .x_out(stage_9_per_in[50]),
    .y_out(stage_9_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_26 (
    .x_in(stage_8_per_out[52]),
    .y_in(stage_8_per_out[53]),
    .x_out(stage_9_per_in[52]),
    .y_out(stage_9_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_27 (
    .x_in(stage_8_per_out[54]),
    .y_in(stage_8_per_out[55]),
    .x_out(stage_9_per_in[54]),
    .y_out(stage_9_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_28 (
    .x_in(stage_8_per_out[56]),
    .y_in(stage_8_per_out[57]),
    .x_out(stage_9_per_in[56]),
    .y_out(stage_9_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_29 (
    .x_in(stage_8_per_out[58]),
    .y_in(stage_8_per_out[59]),
    .x_out(stage_9_per_in[58]),
    .y_out(stage_9_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_30 (
    .x_in(stage_8_per_out[60]),
    .y_in(stage_8_per_out[61]),
    .x_out(stage_9_per_in[60]),
    .y_out(stage_9_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_31 (
    .x_in(stage_8_per_out[62]),
    .y_in(stage_8_per_out[63]),
    .x_out(stage_9_per_in[62]),
    .y_out(stage_9_per_in[63]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_32 (
    .x_in(stage_8_per_out[64]),
    .y_in(stage_8_per_out[65]),
    .x_out(stage_9_per_in[64]),
    .y_out(stage_9_per_in[65]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_33 (
    .x_in(stage_8_per_out[66]),
    .y_in(stage_8_per_out[67]),
    .x_out(stage_9_per_in[66]),
    .y_out(stage_9_per_in[67]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_34 (
    .x_in(stage_8_per_out[68]),
    .y_in(stage_8_per_out[69]),
    .x_out(stage_9_per_in[68]),
    .y_out(stage_9_per_in[69]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_35 (
    .x_in(stage_8_per_out[70]),
    .y_in(stage_8_per_out[71]),
    .x_out(stage_9_per_in[70]),
    .y_out(stage_9_per_in[71]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_36 (
    .x_in(stage_8_per_out[72]),
    .y_in(stage_8_per_out[73]),
    .x_out(stage_9_per_in[72]),
    .y_out(stage_9_per_in[73]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_37 (
    .x_in(stage_8_per_out[74]),
    .y_in(stage_8_per_out[75]),
    .x_out(stage_9_per_in[74]),
    .y_out(stage_9_per_in[75]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_38 (
    .x_in(stage_8_per_out[76]),
    .y_in(stage_8_per_out[77]),
    .x_out(stage_9_per_in[76]),
    .y_out(stage_9_per_in[77]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_39 (
    .x_in(stage_8_per_out[78]),
    .y_in(stage_8_per_out[79]),
    .x_out(stage_9_per_in[78]),
    .y_out(stage_9_per_in[79]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_40 (
    .x_in(stage_8_per_out[80]),
    .y_in(stage_8_per_out[81]),
    .x_out(stage_9_per_in[80]),
    .y_out(stage_9_per_in[81]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_41 (
    .x_in(stage_8_per_out[82]),
    .y_in(stage_8_per_out[83]),
    .x_out(stage_9_per_in[82]),
    .y_out(stage_9_per_in[83]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_42 (
    .x_in(stage_8_per_out[84]),
    .y_in(stage_8_per_out[85]),
    .x_out(stage_9_per_in[84]),
    .y_out(stage_9_per_in[85]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_43 (
    .x_in(stage_8_per_out[86]),
    .y_in(stage_8_per_out[87]),
    .x_out(stage_9_per_in[86]),
    .y_out(stage_9_per_in[87]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_44 (
    .x_in(stage_8_per_out[88]),
    .y_in(stage_8_per_out[89]),
    .x_out(stage_9_per_in[88]),
    .y_out(stage_9_per_in[89]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_45 (
    .x_in(stage_8_per_out[90]),
    .y_in(stage_8_per_out[91]),
    .x_out(stage_9_per_in[90]),
    .y_out(stage_9_per_in[91]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_46 (
    .x_in(stage_8_per_out[92]),
    .y_in(stage_8_per_out[93]),
    .x_out(stage_9_per_in[92]),
    .y_out(stage_9_per_in[93]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_47 (
    .x_in(stage_8_per_out[94]),
    .y_in(stage_8_per_out[95]),
    .x_out(stage_9_per_in[94]),
    .y_out(stage_9_per_in[95]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_48 (
    .x_in(stage_8_per_out[96]),
    .y_in(stage_8_per_out[97]),
    .x_out(stage_9_per_in[96]),
    .y_out(stage_9_per_in[97]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_49 (
    .x_in(stage_8_per_out[98]),
    .y_in(stage_8_per_out[99]),
    .x_out(stage_9_per_in[98]),
    .y_out(stage_9_per_in[99]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_50 (
    .x_in(stage_8_per_out[100]),
    .y_in(stage_8_per_out[101]),
    .x_out(stage_9_per_in[100]),
    .y_out(stage_9_per_in[101]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_51 (
    .x_in(stage_8_per_out[102]),
    .y_in(stage_8_per_out[103]),
    .x_out(stage_9_per_in[102]),
    .y_out(stage_9_per_in[103]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_52 (
    .x_in(stage_8_per_out[104]),
    .y_in(stage_8_per_out[105]),
    .x_out(stage_9_per_in[104]),
    .y_out(stage_9_per_in[105]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_53 (
    .x_in(stage_8_per_out[106]),
    .y_in(stage_8_per_out[107]),
    .x_out(stage_9_per_in[106]),
    .y_out(stage_9_per_in[107]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_54 (
    .x_in(stage_8_per_out[108]),
    .y_in(stage_8_per_out[109]),
    .x_out(stage_9_per_in[108]),
    .y_out(stage_9_per_in[109]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_55 (
    .x_in(stage_8_per_out[110]),
    .y_in(stage_8_per_out[111]),
    .x_out(stage_9_per_in[110]),
    .y_out(stage_9_per_in[111]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_56 (
    .x_in(stage_8_per_out[112]),
    .y_in(stage_8_per_out[113]),
    .x_out(stage_9_per_in[112]),
    .y_out(stage_9_per_in[113]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_57 (
    .x_in(stage_8_per_out[114]),
    .y_in(stage_8_per_out[115]),
    .x_out(stage_9_per_in[114]),
    .y_out(stage_9_per_in[115]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_58 (
    .x_in(stage_8_per_out[116]),
    .y_in(stage_8_per_out[117]),
    .x_out(stage_9_per_in[116]),
    .y_out(stage_9_per_in[117]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_59 (
    .x_in(stage_8_per_out[118]),
    .y_in(stage_8_per_out[119]),
    .x_out(stage_9_per_in[118]),
    .y_out(stage_9_per_in[119]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_60 (
    .x_in(stage_8_per_out[120]),
    .y_in(stage_8_per_out[121]),
    .x_out(stage_9_per_in[120]),
    .y_out(stage_9_per_in[121]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_61 (
    .x_in(stage_8_per_out[122]),
    .y_in(stage_8_per_out[123]),
    .x_out(stage_9_per_in[122]),
    .y_out(stage_9_per_in[123]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_62 (
    .x_in(stage_8_per_out[124]),
    .y_in(stage_8_per_out[125]),
    .x_out(stage_9_per_in[124]),
    .y_out(stage_9_per_in[125]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_63 (
    .x_in(stage_8_per_out[126]),
    .y_in(stage_8_per_out[127]),
    .x_out(stage_9_per_in[126]),
    .y_out(stage_9_per_in[127]),
    .clk(clk),
    .rst(rst)
  );



  // TODO(Yang): stage 8 -> stage 9 permutation
  // FIXME: ignore butterfly units for now.
  stage_9_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_9_10_per (
    .inData_0(stage_9_per_in[0]),
    .inData_1(stage_9_per_in[1]),
    .inData_2(stage_9_per_in[2]),
    .inData_3(stage_9_per_in[3]),
    .inData_4(stage_9_per_in[4]),
    .inData_5(stage_9_per_in[5]),
    .inData_6(stage_9_per_in[6]),
    .inData_7(stage_9_per_in[7]),
    .inData_8(stage_9_per_in[8]),
    .inData_9(stage_9_per_in[9]),
    .inData_10(stage_9_per_in[10]),
    .inData_11(stage_9_per_in[11]),
    .inData_12(stage_9_per_in[12]),
    .inData_13(stage_9_per_in[13]),
    .inData_14(stage_9_per_in[14]),
    .inData_15(stage_9_per_in[15]),
    .inData_16(stage_9_per_in[16]),
    .inData_17(stage_9_per_in[17]),
    .inData_18(stage_9_per_in[18]),
    .inData_19(stage_9_per_in[19]),
    .inData_20(stage_9_per_in[20]),
    .inData_21(stage_9_per_in[21]),
    .inData_22(stage_9_per_in[22]),
    .inData_23(stage_9_per_in[23]),
    .inData_24(stage_9_per_in[24]),
    .inData_25(stage_9_per_in[25]),
    .inData_26(stage_9_per_in[26]),
    .inData_27(stage_9_per_in[27]),
    .inData_28(stage_9_per_in[28]),
    .inData_29(stage_9_per_in[29]),
    .inData_30(stage_9_per_in[30]),
    .inData_31(stage_9_per_in[31]),
    .inData_32(stage_9_per_in[32]),
    .inData_33(stage_9_per_in[33]),
    .inData_34(stage_9_per_in[34]),
    .inData_35(stage_9_per_in[35]),
    .inData_36(stage_9_per_in[36]),
    .inData_37(stage_9_per_in[37]),
    .inData_38(stage_9_per_in[38]),
    .inData_39(stage_9_per_in[39]),
    .inData_40(stage_9_per_in[40]),
    .inData_41(stage_9_per_in[41]),
    .inData_42(stage_9_per_in[42]),
    .inData_43(stage_9_per_in[43]),
    .inData_44(stage_9_per_in[44]),
    .inData_45(stage_9_per_in[45]),
    .inData_46(stage_9_per_in[46]),
    .inData_47(stage_9_per_in[47]),
    .inData_48(stage_9_per_in[48]),
    .inData_49(stage_9_per_in[49]),
    .inData_50(stage_9_per_in[50]),
    .inData_51(stage_9_per_in[51]),
    .inData_52(stage_9_per_in[52]),
    .inData_53(stage_9_per_in[53]),
    .inData_54(stage_9_per_in[54]),
    .inData_55(stage_9_per_in[55]),
    .inData_56(stage_9_per_in[56]),
    .inData_57(stage_9_per_in[57]),
    .inData_58(stage_9_per_in[58]),
    .inData_59(stage_9_per_in[59]),
    .inData_60(stage_9_per_in[60]),
    .inData_61(stage_9_per_in[61]),
    .inData_62(stage_9_per_in[62]),
    .inData_63(stage_9_per_in[63]),
    .inData_64(stage_9_per_in[64]),
    .inData_65(stage_9_per_in[65]),
    .inData_66(stage_9_per_in[66]),
    .inData_67(stage_9_per_in[67]),
    .inData_68(stage_9_per_in[68]),
    .inData_69(stage_9_per_in[69]),
    .inData_70(stage_9_per_in[70]),
    .inData_71(stage_9_per_in[71]),
    .inData_72(stage_9_per_in[72]),
    .inData_73(stage_9_per_in[73]),
    .inData_74(stage_9_per_in[74]),
    .inData_75(stage_9_per_in[75]),
    .inData_76(stage_9_per_in[76]),
    .inData_77(stage_9_per_in[77]),
    .inData_78(stage_9_per_in[78]),
    .inData_79(stage_9_per_in[79]),
    .inData_80(stage_9_per_in[80]),
    .inData_81(stage_9_per_in[81]),
    .inData_82(stage_9_per_in[82]),
    .inData_83(stage_9_per_in[83]),
    .inData_84(stage_9_per_in[84]),
    .inData_85(stage_9_per_in[85]),
    .inData_86(stage_9_per_in[86]),
    .inData_87(stage_9_per_in[87]),
    .inData_88(stage_9_per_in[88]),
    .inData_89(stage_9_per_in[89]),
    .inData_90(stage_9_per_in[90]),
    .inData_91(stage_9_per_in[91]),
    .inData_92(stage_9_per_in[92]),
    .inData_93(stage_9_per_in[93]),
    .inData_94(stage_9_per_in[94]),
    .inData_95(stage_9_per_in[95]),
    .inData_96(stage_9_per_in[96]),
    .inData_97(stage_9_per_in[97]),
    .inData_98(stage_9_per_in[98]),
    .inData_99(stage_9_per_in[99]),
    .inData_100(stage_9_per_in[100]),
    .inData_101(stage_9_per_in[101]),
    .inData_102(stage_9_per_in[102]),
    .inData_103(stage_9_per_in[103]),
    .inData_104(stage_9_per_in[104]),
    .inData_105(stage_9_per_in[105]),
    .inData_106(stage_9_per_in[106]),
    .inData_107(stage_9_per_in[107]),
    .inData_108(stage_9_per_in[108]),
    .inData_109(stage_9_per_in[109]),
    .inData_110(stage_9_per_in[110]),
    .inData_111(stage_9_per_in[111]),
    .inData_112(stage_9_per_in[112]),
    .inData_113(stage_9_per_in[113]),
    .inData_114(stage_9_per_in[114]),
    .inData_115(stage_9_per_in[115]),
    .inData_116(stage_9_per_in[116]),
    .inData_117(stage_9_per_in[117]),
    .inData_118(stage_9_per_in[118]),
    .inData_119(stage_9_per_in[119]),
    .inData_120(stage_9_per_in[120]),
    .inData_121(stage_9_per_in[121]),
    .inData_122(stage_9_per_in[122]),
    .inData_123(stage_9_per_in[123]),
    .inData_124(stage_9_per_in[124]),
    .inData_125(stage_9_per_in[125]),
    .inData_126(stage_9_per_in[126]),
    .inData_127(stage_9_per_in[127]),
    .outData_0(stage_9_per_out[0]),
    .outData_1(stage_9_per_out[1]),
    .outData_2(stage_9_per_out[2]),
    .outData_3(stage_9_per_out[3]),
    .outData_4(stage_9_per_out[4]),
    .outData_5(stage_9_per_out[5]),
    .outData_6(stage_9_per_out[6]),
    .outData_7(stage_9_per_out[7]),
    .outData_8(stage_9_per_out[8]),
    .outData_9(stage_9_per_out[9]),
    .outData_10(stage_9_per_out[10]),
    .outData_11(stage_9_per_out[11]),
    .outData_12(stage_9_per_out[12]),
    .outData_13(stage_9_per_out[13]),
    .outData_14(stage_9_per_out[14]),
    .outData_15(stage_9_per_out[15]),
    .outData_16(stage_9_per_out[16]),
    .outData_17(stage_9_per_out[17]),
    .outData_18(stage_9_per_out[18]),
    .outData_19(stage_9_per_out[19]),
    .outData_20(stage_9_per_out[20]),
    .outData_21(stage_9_per_out[21]),
    .outData_22(stage_9_per_out[22]),
    .outData_23(stage_9_per_out[23]),
    .outData_24(stage_9_per_out[24]),
    .outData_25(stage_9_per_out[25]),
    .outData_26(stage_9_per_out[26]),
    .outData_27(stage_9_per_out[27]),
    .outData_28(stage_9_per_out[28]),
    .outData_29(stage_9_per_out[29]),
    .outData_30(stage_9_per_out[30]),
    .outData_31(stage_9_per_out[31]),
    .outData_32(stage_9_per_out[32]),
    .outData_33(stage_9_per_out[33]),
    .outData_34(stage_9_per_out[34]),
    .outData_35(stage_9_per_out[35]),
    .outData_36(stage_9_per_out[36]),
    .outData_37(stage_9_per_out[37]),
    .outData_38(stage_9_per_out[38]),
    .outData_39(stage_9_per_out[39]),
    .outData_40(stage_9_per_out[40]),
    .outData_41(stage_9_per_out[41]),
    .outData_42(stage_9_per_out[42]),
    .outData_43(stage_9_per_out[43]),
    .outData_44(stage_9_per_out[44]),
    .outData_45(stage_9_per_out[45]),
    .outData_46(stage_9_per_out[46]),
    .outData_47(stage_9_per_out[47]),
    .outData_48(stage_9_per_out[48]),
    .outData_49(stage_9_per_out[49]),
    .outData_50(stage_9_per_out[50]),
    .outData_51(stage_9_per_out[51]),
    .outData_52(stage_9_per_out[52]),
    .outData_53(stage_9_per_out[53]),
    .outData_54(stage_9_per_out[54]),
    .outData_55(stage_9_per_out[55]),
    .outData_56(stage_9_per_out[56]),
    .outData_57(stage_9_per_out[57]),
    .outData_58(stage_9_per_out[58]),
    .outData_59(stage_9_per_out[59]),
    .outData_60(stage_9_per_out[60]),
    .outData_61(stage_9_per_out[61]),
    .outData_62(stage_9_per_out[62]),
    .outData_63(stage_9_per_out[63]),
    .outData_64(stage_9_per_out[64]),
    .outData_65(stage_9_per_out[65]),
    .outData_66(stage_9_per_out[66]),
    .outData_67(stage_9_per_out[67]),
    .outData_68(stage_9_per_out[68]),
    .outData_69(stage_9_per_out[69]),
    .outData_70(stage_9_per_out[70]),
    .outData_71(stage_9_per_out[71]),
    .outData_72(stage_9_per_out[72]),
    .outData_73(stage_9_per_out[73]),
    .outData_74(stage_9_per_out[74]),
    .outData_75(stage_9_per_out[75]),
    .outData_76(stage_9_per_out[76]),
    .outData_77(stage_9_per_out[77]),
    .outData_78(stage_9_per_out[78]),
    .outData_79(stage_9_per_out[79]),
    .outData_80(stage_9_per_out[80]),
    .outData_81(stage_9_per_out[81]),
    .outData_82(stage_9_per_out[82]),
    .outData_83(stage_9_per_out[83]),
    .outData_84(stage_9_per_out[84]),
    .outData_85(stage_9_per_out[85]),
    .outData_86(stage_9_per_out[86]),
    .outData_87(stage_9_per_out[87]),
    .outData_88(stage_9_per_out[88]),
    .outData_89(stage_9_per_out[89]),
    .outData_90(stage_9_per_out[90]),
    .outData_91(stage_9_per_out[91]),
    .outData_92(stage_9_per_out[92]),
    .outData_93(stage_9_per_out[93]),
    .outData_94(stage_9_per_out[94]),
    .outData_95(stage_9_per_out[95]),
    .outData_96(stage_9_per_out[96]),
    .outData_97(stage_9_per_out[97]),
    .outData_98(stage_9_per_out[98]),
    .outData_99(stage_9_per_out[99]),
    .outData_100(stage_9_per_out[100]),
    .outData_101(stage_9_per_out[101]),
    .outData_102(stage_9_per_out[102]),
    .outData_103(stage_9_per_out[103]),
    .outData_104(stage_9_per_out[104]),
    .outData_105(stage_9_per_out[105]),
    .outData_106(stage_9_per_out[106]),
    .outData_107(stage_9_per_out[107]),
    .outData_108(stage_9_per_out[108]),
    .outData_109(stage_9_per_out[109]),
    .outData_110(stage_9_per_out[110]),
    .outData_111(stage_9_per_out[111]),
    .outData_112(stage_9_per_out[112]),
    .outData_113(stage_9_per_out[113]),
    .outData_114(stage_9_per_out[114]),
    .outData_115(stage_9_per_out[115]),
    .outData_116(stage_9_per_out[116]),
    .outData_117(stage_9_per_out[117]),
    .outData_118(stage_9_per_out[118]),
    .outData_119(stage_9_per_out[119]),
    .outData_120(stage_9_per_out[120]),
    .outData_121(stage_9_per_out[121]),
    .outData_122(stage_9_per_out[122]),
    .outData_123(stage_9_per_out[123]),
    .outData_124(stage_9_per_out[124]),
    .outData_125(stage_9_per_out[125]),
    .outData_126(stage_9_per_out[126]),
    .outData_127(stage_9_per_out[127]),
    .in_start(in_start[9]),
    .out_start(out_start[9]),
    .clk(clk),
    .rst(rst)
  );

  // TODO(Tian): stage 9 32 butterfly units
  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_0 (
    .x_in(stage_9_per_out[0]),
    .y_in(stage_9_per_out[1]),
    .x_out(stage_10_per_in[0]),
    .y_out(stage_10_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_1 (
    .x_in(stage_9_per_out[2]),
    .y_in(stage_9_per_out[3]),
    .x_out(stage_10_per_in[2]),
    .y_out(stage_10_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_2 (
    .x_in(stage_9_per_out[4]),
    .y_in(stage_9_per_out[5]),
    .x_out(stage_10_per_in[4]),
    .y_out(stage_10_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_3 (
    .x_in(stage_9_per_out[6]),
    .y_in(stage_9_per_out[7]),
    .x_out(stage_10_per_in[6]),
    .y_out(stage_10_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_4 (
    .x_in(stage_9_per_out[8]),
    .y_in(stage_9_per_out[9]),
    .x_out(stage_10_per_in[8]),
    .y_out(stage_10_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_5 (
    .x_in(stage_9_per_out[10]),
    .y_in(stage_9_per_out[11]),
    .x_out(stage_10_per_in[10]),
    .y_out(stage_10_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_6 (
    .x_in(stage_9_per_out[12]),
    .y_in(stage_9_per_out[13]),
    .x_out(stage_10_per_in[12]),
    .y_out(stage_10_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_7 (
    .x_in(stage_9_per_out[14]),
    .y_in(stage_9_per_out[15]),
    .x_out(stage_10_per_in[14]),
    .y_out(stage_10_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_8 (
    .x_in(stage_9_per_out[16]),
    .y_in(stage_9_per_out[17]),
    .x_out(stage_10_per_in[16]),
    .y_out(stage_10_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_9 (
    .x_in(stage_9_per_out[18]),
    .y_in(stage_9_per_out[19]),
    .x_out(stage_10_per_in[18]),
    .y_out(stage_10_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_10 (
    .x_in(stage_9_per_out[20]),
    .y_in(stage_9_per_out[21]),
    .x_out(stage_10_per_in[20]),
    .y_out(stage_10_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_11 (
    .x_in(stage_9_per_out[22]),
    .y_in(stage_9_per_out[23]),
    .x_out(stage_10_per_in[22]),
    .y_out(stage_10_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_12 (
    .x_in(stage_9_per_out[24]),
    .y_in(stage_9_per_out[25]),
    .x_out(stage_10_per_in[24]),
    .y_out(stage_10_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_13 (
    .x_in(stage_9_per_out[26]),
    .y_in(stage_9_per_out[27]),
    .x_out(stage_10_per_in[26]),
    .y_out(stage_10_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_14 (
    .x_in(stage_9_per_out[28]),
    .y_in(stage_9_per_out[29]),
    .x_out(stage_10_per_in[28]),
    .y_out(stage_10_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_15 (
    .x_in(stage_9_per_out[30]),
    .y_in(stage_9_per_out[31]),
    .x_out(stage_10_per_in[30]),
    .y_out(stage_10_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_16 (
    .x_in(stage_9_per_out[32]),
    .y_in(stage_9_per_out[33]),
    .x_out(stage_10_per_in[32]),
    .y_out(stage_10_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_17 (
    .x_in(stage_9_per_out[34]),
    .y_in(stage_9_per_out[35]),
    .x_out(stage_10_per_in[34]),
    .y_out(stage_10_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_18 (
    .x_in(stage_9_per_out[36]),
    .y_in(stage_9_per_out[37]),
    .x_out(stage_10_per_in[36]),
    .y_out(stage_10_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_19 (
    .x_in(stage_9_per_out[38]),
    .y_in(stage_9_per_out[39]),
    .x_out(stage_10_per_in[38]),
    .y_out(stage_10_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_20 (
    .x_in(stage_9_per_out[40]),
    .y_in(stage_9_per_out[41]),
    .x_out(stage_10_per_in[40]),
    .y_out(stage_10_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_21 (
    .x_in(stage_9_per_out[42]),
    .y_in(stage_9_per_out[43]),
    .x_out(stage_10_per_in[42]),
    .y_out(stage_10_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_22 (
    .x_in(stage_9_per_out[44]),
    .y_in(stage_9_per_out[45]),
    .x_out(stage_10_per_in[44]),
    .y_out(stage_10_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_23 (
    .x_in(stage_9_per_out[46]),
    .y_in(stage_9_per_out[47]),
    .x_out(stage_10_per_in[46]),
    .y_out(stage_10_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_24 (
    .x_in(stage_9_per_out[48]),
    .y_in(stage_9_per_out[49]),
    .x_out(stage_10_per_in[48]),
    .y_out(stage_10_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_25 (
    .x_in(stage_9_per_out[50]),
    .y_in(stage_9_per_out[51]),
    .x_out(stage_10_per_in[50]),
    .y_out(stage_10_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_26 (
    .x_in(stage_9_per_out[52]),
    .y_in(stage_9_per_out[53]),
    .x_out(stage_10_per_in[52]),
    .y_out(stage_10_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_27 (
    .x_in(stage_9_per_out[54]),
    .y_in(stage_9_per_out[55]),
    .x_out(stage_10_per_in[54]),
    .y_out(stage_10_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_28 (
    .x_in(stage_9_per_out[56]),
    .y_in(stage_9_per_out[57]),
    .x_out(stage_10_per_in[56]),
    .y_out(stage_10_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_29 (
    .x_in(stage_9_per_out[58]),
    .y_in(stage_9_per_out[59]),
    .x_out(stage_10_per_in[58]),
    .y_out(stage_10_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_30 (
    .x_in(stage_9_per_out[60]),
    .y_in(stage_9_per_out[61]),
    .x_out(stage_10_per_in[60]),
    .y_out(stage_10_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_31 (
    .x_in(stage_9_per_out[62]),
    .y_in(stage_9_per_out[63]),
    .x_out(stage_10_per_in[62]),
    .y_out(stage_10_per_in[63]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_32 (
    .x_in(stage_9_per_out[64]),
    .y_in(stage_9_per_out[65]),
    .x_out(stage_10_per_in[64]),
    .y_out(stage_10_per_in[65]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_33 (
    .x_in(stage_9_per_out[66]),
    .y_in(stage_9_per_out[67]),
    .x_out(stage_10_per_in[66]),
    .y_out(stage_10_per_in[67]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_34 (
    .x_in(stage_9_per_out[68]),
    .y_in(stage_9_per_out[69]),
    .x_out(stage_10_per_in[68]),
    .y_out(stage_10_per_in[69]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_35 (
    .x_in(stage_9_per_out[70]),
    .y_in(stage_9_per_out[71]),
    .x_out(stage_10_per_in[70]),
    .y_out(stage_10_per_in[71]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_36 (
    .x_in(stage_9_per_out[72]),
    .y_in(stage_9_per_out[73]),
    .x_out(stage_10_per_in[72]),
    .y_out(stage_10_per_in[73]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_37 (
    .x_in(stage_9_per_out[74]),
    .y_in(stage_9_per_out[75]),
    .x_out(stage_10_per_in[74]),
    .y_out(stage_10_per_in[75]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_38 (
    .x_in(stage_9_per_out[76]),
    .y_in(stage_9_per_out[77]),
    .x_out(stage_10_per_in[76]),
    .y_out(stage_10_per_in[77]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_39 (
    .x_in(stage_9_per_out[78]),
    .y_in(stage_9_per_out[79]),
    .x_out(stage_10_per_in[78]),
    .y_out(stage_10_per_in[79]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_40 (
    .x_in(stage_9_per_out[80]),
    .y_in(stage_9_per_out[81]),
    .x_out(stage_10_per_in[80]),
    .y_out(stage_10_per_in[81]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_41 (
    .x_in(stage_9_per_out[82]),
    .y_in(stage_9_per_out[83]),
    .x_out(stage_10_per_in[82]),
    .y_out(stage_10_per_in[83]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_42 (
    .x_in(stage_9_per_out[84]),
    .y_in(stage_9_per_out[85]),
    .x_out(stage_10_per_in[84]),
    .y_out(stage_10_per_in[85]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_43 (
    .x_in(stage_9_per_out[86]),
    .y_in(stage_9_per_out[87]),
    .x_out(stage_10_per_in[86]),
    .y_out(stage_10_per_in[87]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_44 (
    .x_in(stage_9_per_out[88]),
    .y_in(stage_9_per_out[89]),
    .x_out(stage_10_per_in[88]),
    .y_out(stage_10_per_in[89]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_45 (
    .x_in(stage_9_per_out[90]),
    .y_in(stage_9_per_out[91]),
    .x_out(stage_10_per_in[90]),
    .y_out(stage_10_per_in[91]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_46 (
    .x_in(stage_9_per_out[92]),
    .y_in(stage_9_per_out[93]),
    .x_out(stage_10_per_in[92]),
    .y_out(stage_10_per_in[93]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_47 (
    .x_in(stage_9_per_out[94]),
    .y_in(stage_9_per_out[95]),
    .x_out(stage_10_per_in[94]),
    .y_out(stage_10_per_in[95]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_48 (
    .x_in(stage_9_per_out[96]),
    .y_in(stage_9_per_out[97]),
    .x_out(stage_10_per_in[96]),
    .y_out(stage_10_per_in[97]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_49 (
    .x_in(stage_9_per_out[98]),
    .y_in(stage_9_per_out[99]),
    .x_out(stage_10_per_in[98]),
    .y_out(stage_10_per_in[99]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_50 (
    .x_in(stage_9_per_out[100]),
    .y_in(stage_9_per_out[101]),
    .x_out(stage_10_per_in[100]),
    .y_out(stage_10_per_in[101]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_51 (
    .x_in(stage_9_per_out[102]),
    .y_in(stage_9_per_out[103]),
    .x_out(stage_10_per_in[102]),
    .y_out(stage_10_per_in[103]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_52 (
    .x_in(stage_9_per_out[104]),
    .y_in(stage_9_per_out[105]),
    .x_out(stage_10_per_in[104]),
    .y_out(stage_10_per_in[105]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_53 (
    .x_in(stage_9_per_out[106]),
    .y_in(stage_9_per_out[107]),
    .x_out(stage_10_per_in[106]),
    .y_out(stage_10_per_in[107]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_54 (
    .x_in(stage_9_per_out[108]),
    .y_in(stage_9_per_out[109]),
    .x_out(stage_10_per_in[108]),
    .y_out(stage_10_per_in[109]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_55 (
    .x_in(stage_9_per_out[110]),
    .y_in(stage_9_per_out[111]),
    .x_out(stage_10_per_in[110]),
    .y_out(stage_10_per_in[111]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_56 (
    .x_in(stage_9_per_out[112]),
    .y_in(stage_9_per_out[113]),
    .x_out(stage_10_per_in[112]),
    .y_out(stage_10_per_in[113]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_57 (
    .x_in(stage_9_per_out[114]),
    .y_in(stage_9_per_out[115]),
    .x_out(stage_10_per_in[114]),
    .y_out(stage_10_per_in[115]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_58 (
    .x_in(stage_9_per_out[116]),
    .y_in(stage_9_per_out[117]),
    .x_out(stage_10_per_in[116]),
    .y_out(stage_10_per_in[117]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_59 (
    .x_in(stage_9_per_out[118]),
    .y_in(stage_9_per_out[119]),
    .x_out(stage_10_per_in[118]),
    .y_out(stage_10_per_in[119]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_60 (
    .x_in(stage_9_per_out[120]),
    .y_in(stage_9_per_out[121]),
    .x_out(stage_10_per_in[120]),
    .y_out(stage_10_per_in[121]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_61 (
    .x_in(stage_9_per_out[122]),
    .y_in(stage_9_per_out[123]),
    .x_out(stage_10_per_in[122]),
    .y_out(stage_10_per_in[123]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_62 (
    .x_in(stage_9_per_out[124]),
    .y_in(stage_9_per_out[125]),
    .x_out(stage_10_per_in[124]),
    .y_out(stage_10_per_in[125]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_63 (
    .x_in(stage_9_per_out[126]),
    .y_in(stage_9_per_out[127]),
    .x_out(stage_10_per_in[126]),
    .y_out(stage_10_per_in[127]),
    .clk(clk),
    .rst(rst)
  );



  // TODO(Yang): stage 8 -> stage 9 permutation
  // FIXME: ignore butterfly units for now.
  stage_10_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_10_11_per (
    .inData_0(stage_10_per_in[0]),
    .inData_1(stage_10_per_in[1]),
    .inData_2(stage_10_per_in[2]),
    .inData_3(stage_10_per_in[3]),
    .inData_4(stage_10_per_in[4]),
    .inData_5(stage_10_per_in[5]),
    .inData_6(stage_10_per_in[6]),
    .inData_7(stage_10_per_in[7]),
    .inData_8(stage_10_per_in[8]),
    .inData_9(stage_10_per_in[9]),
    .inData_10(stage_10_per_in[10]),
    .inData_11(stage_10_per_in[11]),
    .inData_12(stage_10_per_in[12]),
    .inData_13(stage_10_per_in[13]),
    .inData_14(stage_10_per_in[14]),
    .inData_15(stage_10_per_in[15]),
    .inData_16(stage_10_per_in[16]),
    .inData_17(stage_10_per_in[17]),
    .inData_18(stage_10_per_in[18]),
    .inData_19(stage_10_per_in[19]),
    .inData_20(stage_10_per_in[20]),
    .inData_21(stage_10_per_in[21]),
    .inData_22(stage_10_per_in[22]),
    .inData_23(stage_10_per_in[23]),
    .inData_24(stage_10_per_in[24]),
    .inData_25(stage_10_per_in[25]),
    .inData_26(stage_10_per_in[26]),
    .inData_27(stage_10_per_in[27]),
    .inData_28(stage_10_per_in[28]),
    .inData_29(stage_10_per_in[29]),
    .inData_30(stage_10_per_in[30]),
    .inData_31(stage_10_per_in[31]),
    .inData_32(stage_10_per_in[32]),
    .inData_33(stage_10_per_in[33]),
    .inData_34(stage_10_per_in[34]),
    .inData_35(stage_10_per_in[35]),
    .inData_36(stage_10_per_in[36]),
    .inData_37(stage_10_per_in[37]),
    .inData_38(stage_10_per_in[38]),
    .inData_39(stage_10_per_in[39]),
    .inData_40(stage_10_per_in[40]),
    .inData_41(stage_10_per_in[41]),
    .inData_42(stage_10_per_in[42]),
    .inData_43(stage_10_per_in[43]),
    .inData_44(stage_10_per_in[44]),
    .inData_45(stage_10_per_in[45]),
    .inData_46(stage_10_per_in[46]),
    .inData_47(stage_10_per_in[47]),
    .inData_48(stage_10_per_in[48]),
    .inData_49(stage_10_per_in[49]),
    .inData_50(stage_10_per_in[50]),
    .inData_51(stage_10_per_in[51]),
    .inData_52(stage_10_per_in[52]),
    .inData_53(stage_10_per_in[53]),
    .inData_54(stage_10_per_in[54]),
    .inData_55(stage_10_per_in[55]),
    .inData_56(stage_10_per_in[56]),
    .inData_57(stage_10_per_in[57]),
    .inData_58(stage_10_per_in[58]),
    .inData_59(stage_10_per_in[59]),
    .inData_60(stage_10_per_in[60]),
    .inData_61(stage_10_per_in[61]),
    .inData_62(stage_10_per_in[62]),
    .inData_63(stage_10_per_in[63]),
    .inData_64(stage_10_per_in[64]),
    .inData_65(stage_10_per_in[65]),
    .inData_66(stage_10_per_in[66]),
    .inData_67(stage_10_per_in[67]),
    .inData_68(stage_10_per_in[68]),
    .inData_69(stage_10_per_in[69]),
    .inData_70(stage_10_per_in[70]),
    .inData_71(stage_10_per_in[71]),
    .inData_72(stage_10_per_in[72]),
    .inData_73(stage_10_per_in[73]),
    .inData_74(stage_10_per_in[74]),
    .inData_75(stage_10_per_in[75]),
    .inData_76(stage_10_per_in[76]),
    .inData_77(stage_10_per_in[77]),
    .inData_78(stage_10_per_in[78]),
    .inData_79(stage_10_per_in[79]),
    .inData_80(stage_10_per_in[80]),
    .inData_81(stage_10_per_in[81]),
    .inData_82(stage_10_per_in[82]),
    .inData_83(stage_10_per_in[83]),
    .inData_84(stage_10_per_in[84]),
    .inData_85(stage_10_per_in[85]),
    .inData_86(stage_10_per_in[86]),
    .inData_87(stage_10_per_in[87]),
    .inData_88(stage_10_per_in[88]),
    .inData_89(stage_10_per_in[89]),
    .inData_90(stage_10_per_in[90]),
    .inData_91(stage_10_per_in[91]),
    .inData_92(stage_10_per_in[92]),
    .inData_93(stage_10_per_in[93]),
    .inData_94(stage_10_per_in[94]),
    .inData_95(stage_10_per_in[95]),
    .inData_96(stage_10_per_in[96]),
    .inData_97(stage_10_per_in[97]),
    .inData_98(stage_10_per_in[98]),
    .inData_99(stage_10_per_in[99]),
    .inData_100(stage_10_per_in[100]),
    .inData_101(stage_10_per_in[101]),
    .inData_102(stage_10_per_in[102]),
    .inData_103(stage_10_per_in[103]),
    .inData_104(stage_10_per_in[104]),
    .inData_105(stage_10_per_in[105]),
    .inData_106(stage_10_per_in[106]),
    .inData_107(stage_10_per_in[107]),
    .inData_108(stage_10_per_in[108]),
    .inData_109(stage_10_per_in[109]),
    .inData_110(stage_10_per_in[110]),
    .inData_111(stage_10_per_in[111]),
    .inData_112(stage_10_per_in[112]),
    .inData_113(stage_10_per_in[113]),
    .inData_114(stage_10_per_in[114]),
    .inData_115(stage_10_per_in[115]),
    .inData_116(stage_10_per_in[116]),
    .inData_117(stage_10_per_in[117]),
    .inData_118(stage_10_per_in[118]),
    .inData_119(stage_10_per_in[119]),
    .inData_120(stage_10_per_in[120]),
    .inData_121(stage_10_per_in[121]),
    .inData_122(stage_10_per_in[122]),
    .inData_123(stage_10_per_in[123]),
    .inData_124(stage_10_per_in[124]),
    .inData_125(stage_10_per_in[125]),
    .inData_126(stage_10_per_in[126]),
    .inData_127(stage_10_per_in[127]),
    .outData_0(stage_10_per_out[0]),
    .outData_1(stage_10_per_out[1]),
    .outData_2(stage_10_per_out[2]),
    .outData_3(stage_10_per_out[3]),
    .outData_4(stage_10_per_out[4]),
    .outData_5(stage_10_per_out[5]),
    .outData_6(stage_10_per_out[6]),
    .outData_7(stage_10_per_out[7]),
    .outData_8(stage_10_per_out[8]),
    .outData_9(stage_10_per_out[9]),
    .outData_10(stage_10_per_out[10]),
    .outData_11(stage_10_per_out[11]),
    .outData_12(stage_10_per_out[12]),
    .outData_13(stage_10_per_out[13]),
    .outData_14(stage_10_per_out[14]),
    .outData_15(stage_10_per_out[15]),
    .outData_16(stage_10_per_out[16]),
    .outData_17(stage_10_per_out[17]),
    .outData_18(stage_10_per_out[18]),
    .outData_19(stage_10_per_out[19]),
    .outData_20(stage_10_per_out[20]),
    .outData_21(stage_10_per_out[21]),
    .outData_22(stage_10_per_out[22]),
    .outData_23(stage_10_per_out[23]),
    .outData_24(stage_10_per_out[24]),
    .outData_25(stage_10_per_out[25]),
    .outData_26(stage_10_per_out[26]),
    .outData_27(stage_10_per_out[27]),
    .outData_28(stage_10_per_out[28]),
    .outData_29(stage_10_per_out[29]),
    .outData_30(stage_10_per_out[30]),
    .outData_31(stage_10_per_out[31]),
    .outData_32(stage_10_per_out[32]),
    .outData_33(stage_10_per_out[33]),
    .outData_34(stage_10_per_out[34]),
    .outData_35(stage_10_per_out[35]),
    .outData_36(stage_10_per_out[36]),
    .outData_37(stage_10_per_out[37]),
    .outData_38(stage_10_per_out[38]),
    .outData_39(stage_10_per_out[39]),
    .outData_40(stage_10_per_out[40]),
    .outData_41(stage_10_per_out[41]),
    .outData_42(stage_10_per_out[42]),
    .outData_43(stage_10_per_out[43]),
    .outData_44(stage_10_per_out[44]),
    .outData_45(stage_10_per_out[45]),
    .outData_46(stage_10_per_out[46]),
    .outData_47(stage_10_per_out[47]),
    .outData_48(stage_10_per_out[48]),
    .outData_49(stage_10_per_out[49]),
    .outData_50(stage_10_per_out[50]),
    .outData_51(stage_10_per_out[51]),
    .outData_52(stage_10_per_out[52]),
    .outData_53(stage_10_per_out[53]),
    .outData_54(stage_10_per_out[54]),
    .outData_55(stage_10_per_out[55]),
    .outData_56(stage_10_per_out[56]),
    .outData_57(stage_10_per_out[57]),
    .outData_58(stage_10_per_out[58]),
    .outData_59(stage_10_per_out[59]),
    .outData_60(stage_10_per_out[60]),
    .outData_61(stage_10_per_out[61]),
    .outData_62(stage_10_per_out[62]),
    .outData_63(stage_10_per_out[63]),
    .outData_64(stage_10_per_out[64]),
    .outData_65(stage_10_per_out[65]),
    .outData_66(stage_10_per_out[66]),
    .outData_67(stage_10_per_out[67]),
    .outData_68(stage_10_per_out[68]),
    .outData_69(stage_10_per_out[69]),
    .outData_70(stage_10_per_out[70]),
    .outData_71(stage_10_per_out[71]),
    .outData_72(stage_10_per_out[72]),
    .outData_73(stage_10_per_out[73]),
    .outData_74(stage_10_per_out[74]),
    .outData_75(stage_10_per_out[75]),
    .outData_76(stage_10_per_out[76]),
    .outData_77(stage_10_per_out[77]),
    .outData_78(stage_10_per_out[78]),
    .outData_79(stage_10_per_out[79]),
    .outData_80(stage_10_per_out[80]),
    .outData_81(stage_10_per_out[81]),
    .outData_82(stage_10_per_out[82]),
    .outData_83(stage_10_per_out[83]),
    .outData_84(stage_10_per_out[84]),
    .outData_85(stage_10_per_out[85]),
    .outData_86(stage_10_per_out[86]),
    .outData_87(stage_10_per_out[87]),
    .outData_88(stage_10_per_out[88]),
    .outData_89(stage_10_per_out[89]),
    .outData_90(stage_10_per_out[90]),
    .outData_91(stage_10_per_out[91]),
    .outData_92(stage_10_per_out[92]),
    .outData_93(stage_10_per_out[93]),
    .outData_94(stage_10_per_out[94]),
    .outData_95(stage_10_per_out[95]),
    .outData_96(stage_10_per_out[96]),
    .outData_97(stage_10_per_out[97]),
    .outData_98(stage_10_per_out[98]),
    .outData_99(stage_10_per_out[99]),
    .outData_100(stage_10_per_out[100]),
    .outData_101(stage_10_per_out[101]),
    .outData_102(stage_10_per_out[102]),
    .outData_103(stage_10_per_out[103]),
    .outData_104(stage_10_per_out[104]),
    .outData_105(stage_10_per_out[105]),
    .outData_106(stage_10_per_out[106]),
    .outData_107(stage_10_per_out[107]),
    .outData_108(stage_10_per_out[108]),
    .outData_109(stage_10_per_out[109]),
    .outData_110(stage_10_per_out[110]),
    .outData_111(stage_10_per_out[111]),
    .outData_112(stage_10_per_out[112]),
    .outData_113(stage_10_per_out[113]),
    .outData_114(stage_10_per_out[114]),
    .outData_115(stage_10_per_out[115]),
    .outData_116(stage_10_per_out[116]),
    .outData_117(stage_10_per_out[117]),
    .outData_118(stage_10_per_out[118]),
    .outData_119(stage_10_per_out[119]),
    .outData_120(stage_10_per_out[120]),
    .outData_121(stage_10_per_out[121]),
    .outData_122(stage_10_per_out[122]),
    .outData_123(stage_10_per_out[123]),
    .outData_124(stage_10_per_out[124]),
    .outData_125(stage_10_per_out[125]),
    .outData_126(stage_10_per_out[126]),
    .outData_127(stage_10_per_out[127]),
    .in_start(in_start[10]),
    .out_start(out_start[10]),
    .clk(clk),
    .rst(rst)
  );

  // TODO(Tian): stage 9 32 butterfly units
  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_0 (
    .x_in(stage_10_per_out[0]),
    .y_in(stage_10_per_out[1]),
    .x_out(outData[0]),
    .y_out(outData[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_1 (
    .x_in(stage_10_per_out[2]),
    .y_in(stage_10_per_out[3]),
    .x_out(outData[2]),
    .y_out(outData[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_2 (
    .x_in(stage_10_per_out[4]),
    .y_in(stage_10_per_out[5]),
    .x_out(outData[4]),
    .y_out(outData[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_3 (
    .x_in(stage_10_per_out[6]),
    .y_in(stage_10_per_out[7]),
    .x_out(outData[6]),
    .y_out(outData[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_4 (
    .x_in(stage_10_per_out[8]),
    .y_in(stage_10_per_out[9]),
    .x_out(outData[8]),
    .y_out(outData[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_5 (
    .x_in(stage_10_per_out[10]),
    .y_in(stage_10_per_out[11]),
    .x_out(outData[10]),
    .y_out(outData[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_6 (
    .x_in(stage_10_per_out[12]),
    .y_in(stage_10_per_out[13]),
    .x_out(outData[12]),
    .y_out(outData[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_7 (
    .x_in(stage_10_per_out[14]),
    .y_in(stage_10_per_out[15]),
    .x_out(outData[14]),
    .y_out(outData[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_8 (
    .x_in(stage_10_per_out[16]),
    .y_in(stage_10_per_out[17]),
    .x_out(outData[16]),
    .y_out(outData[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_9 (
    .x_in(stage_10_per_out[18]),
    .y_in(stage_10_per_out[19]),
    .x_out(outData[18]),
    .y_out(outData[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_10 (
    .x_in(stage_10_per_out[20]),
    .y_in(stage_10_per_out[21]),
    .x_out(outData[20]),
    .y_out(outData[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_11 (
    .x_in(stage_10_per_out[22]),
    .y_in(stage_10_per_out[23]),
    .x_out(outData[22]),
    .y_out(outData[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_12 (
    .x_in(stage_10_per_out[24]),
    .y_in(stage_10_per_out[25]),
    .x_out(outData[24]),
    .y_out(outData[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_13 (
    .x_in(stage_10_per_out[26]),
    .y_in(stage_10_per_out[27]),
    .x_out(outData[26]),
    .y_out(outData[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_14 (
    .x_in(stage_10_per_out[28]),
    .y_in(stage_10_per_out[29]),
    .x_out(outData[28]),
    .y_out(outData[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_15 (
    .x_in(stage_10_per_out[30]),
    .y_in(stage_10_per_out[31]),
    .x_out(outData[30]),
    .y_out(outData[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_16 (
    .x_in(stage_10_per_out[32]),
    .y_in(stage_10_per_out[33]),
    .x_out(outData[32]),
    .y_out(outData[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_17 (
    .x_in(stage_10_per_out[34]),
    .y_in(stage_10_per_out[35]),
    .x_out(outData[34]),
    .y_out(outData[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_18 (
    .x_in(stage_10_per_out[36]),
    .y_in(stage_10_per_out[37]),
    .x_out(outData[36]),
    .y_out(outData[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_19 (
    .x_in(stage_10_per_out[38]),
    .y_in(stage_10_per_out[39]),
    .x_out(outData[38]),
    .y_out(outData[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_20 (
    .x_in(stage_10_per_out[40]),
    .y_in(stage_10_per_out[41]),
    .x_out(outData[40]),
    .y_out(outData[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_21 (
    .x_in(stage_10_per_out[42]),
    .y_in(stage_10_per_out[43]),
    .x_out(outData[42]),
    .y_out(outData[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_22 (
    .x_in(stage_10_per_out[44]),
    .y_in(stage_10_per_out[45]),
    .x_out(outData[44]),
    .y_out(outData[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_23 (
    .x_in(stage_10_per_out[46]),
    .y_in(stage_10_per_out[47]),
    .x_out(outData[46]),
    .y_out(outData[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_24 (
    .x_in(stage_10_per_out[48]),
    .y_in(stage_10_per_out[49]),
    .x_out(outData[48]),
    .y_out(outData[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_25 (
    .x_in(stage_10_per_out[50]),
    .y_in(stage_10_per_out[51]),
    .x_out(outData[50]),
    .y_out(outData[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_26 (
    .x_in(stage_10_per_out[52]),
    .y_in(stage_10_per_out[53]),
    .x_out(outData[52]),
    .y_out(outData[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_27 (
    .x_in(stage_10_per_out[54]),
    .y_in(stage_10_per_out[55]),
    .x_out(outData[54]),
    .y_out(outData[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_28 (
    .x_in(stage_10_per_out[56]),
    .y_in(stage_10_per_out[57]),
    .x_out(outData[56]),
    .y_out(outData[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_29 (
    .x_in(stage_10_per_out[58]),
    .y_in(stage_10_per_out[59]),
    .x_out(outData[58]),
    .y_out(outData[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_30 (
    .x_in(stage_10_per_out[60]),
    .y_in(stage_10_per_out[61]),
    .x_out(outData[60]),
    .y_out(outData[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_31 (
    .x_in(stage_10_per_out[62]),
    .y_in(stage_10_per_out[63]),
    .x_out(outData[62]),
    .y_out(outData[63]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_32 (
    .x_in(stage_10_per_out[64]),
    .y_in(stage_10_per_out[65]),
    .x_out(outData[64]),
    .y_out(outData[65]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_33 (
    .x_in(stage_10_per_out[66]),
    .y_in(stage_10_per_out[67]),
    .x_out(outData[66]),
    .y_out(outData[67]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_34 (
    .x_in(stage_10_per_out[68]),
    .y_in(stage_10_per_out[69]),
    .x_out(outData[68]),
    .y_out(outData[69]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_35 (
    .x_in(stage_10_per_out[70]),
    .y_in(stage_10_per_out[71]),
    .x_out(outData[70]),
    .y_out(outData[71]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_36 (
    .x_in(stage_10_per_out[72]),
    .y_in(stage_10_per_out[73]),
    .x_out(outData[72]),
    .y_out(outData[73]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_37 (
    .x_in(stage_10_per_out[74]),
    .y_in(stage_10_per_out[75]),
    .x_out(outData[74]),
    .y_out(outData[75]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_38 (
    .x_in(stage_10_per_out[76]),
    .y_in(stage_10_per_out[77]),
    .x_out(outData[76]),
    .y_out(outData[77]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_39 (
    .x_in(stage_10_per_out[78]),
    .y_in(stage_10_per_out[79]),
    .x_out(outData[78]),
    .y_out(outData[79]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_40 (
    .x_in(stage_10_per_out[80]),
    .y_in(stage_10_per_out[81]),
    .x_out(outData[80]),
    .y_out(outData[81]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_41 (
    .x_in(stage_10_per_out[82]),
    .y_in(stage_10_per_out[83]),
    .x_out(outData[82]),
    .y_out(outData[83]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_42 (
    .x_in(stage_10_per_out[84]),
    .y_in(stage_10_per_out[85]),
    .x_out(outData[84]),
    .y_out(outData[85]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_43 (
    .x_in(stage_10_per_out[86]),
    .y_in(stage_10_per_out[87]),
    .x_out(outData[86]),
    .y_out(outData[87]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_44 (
    .x_in(stage_10_per_out[88]),
    .y_in(stage_10_per_out[89]),
    .x_out(outData[88]),
    .y_out(outData[89]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_45 (
    .x_in(stage_10_per_out[90]),
    .y_in(stage_10_per_out[91]),
    .x_out(outData[90]),
    .y_out(outData[91]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_46 (
    .x_in(stage_10_per_out[92]),
    .y_in(stage_10_per_out[93]),
    .x_out(outData[92]),
    .y_out(outData[93]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_47 (
    .x_in(stage_10_per_out[94]),
    .y_in(stage_10_per_out[95]),
    .x_out(outData[94]),
    .y_out(outData[95]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_48 (
    .x_in(stage_10_per_out[96]),
    .y_in(stage_10_per_out[97]),
    .x_out(outData[96]),
    .y_out(outData[97]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_49 (
    .x_in(stage_10_per_out[98]),
    .y_in(stage_10_per_out[99]),
    .x_out(outData[98]),
    .y_out(outData[99]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_50 (
    .x_in(stage_10_per_out[100]),
    .y_in(stage_10_per_out[101]),
    .x_out(outData[100]),
    .y_out(outData[101]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_51 (
    .x_in(stage_10_per_out[102]),
    .y_in(stage_10_per_out[103]),
    .x_out(outData[102]),
    .y_out(outData[103]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_52 (
    .x_in(stage_10_per_out[104]),
    .y_in(stage_10_per_out[105]),
    .x_out(outData[104]),
    .y_out(outData[105]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_53 (
    .x_in(stage_10_per_out[106]),
    .y_in(stage_10_per_out[107]),
    .x_out(outData[106]),
    .y_out(outData[107]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_54 (
    .x_in(stage_10_per_out[108]),
    .y_in(stage_10_per_out[109]),
    .x_out(outData[108]),
    .y_out(outData[109]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_55 (
    .x_in(stage_10_per_out[110]),
    .y_in(stage_10_per_out[111]),
    .x_out(outData[110]),
    .y_out(outData[111]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_56 (
    .x_in(stage_10_per_out[112]),
    .y_in(stage_10_per_out[113]),
    .x_out(outData[112]),
    .y_out(outData[113]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_57 (
    .x_in(stage_10_per_out[114]),
    .y_in(stage_10_per_out[115]),
    .x_out(outData[114]),
    .y_out(outData[115]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_58 (
    .x_in(stage_10_per_out[116]),
    .y_in(stage_10_per_out[117]),
    .x_out(outData[116]),
    .y_out(outData[117]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_59 (
    .x_in(stage_10_per_out[118]),
    .y_in(stage_10_per_out[119]),
    .x_out(outData[118]),
    .y_out(outData[119]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_60 (
    .x_in(stage_10_per_out[120]),
    .y_in(stage_10_per_out[121]),
    .x_out(outData[120]),
    .y_out(outData[121]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_61 (
    .x_in(stage_10_per_out[122]),
    .y_in(stage_10_per_out[123]),
    .x_out(outData[122]),
    .y_out(outData[123]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_62 (
    .x_in(stage_10_per_out[124]),
    .y_in(stage_10_per_out[125]),
    .x_out(outData[124]),
    .y_out(outData[125]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_63 (
    .x_in(stage_10_per_out[126]),
    .y_in(stage_10_per_out[127]),
    .x_out(outData[126]),
    .y_out(outData[127]),
    .clk(clk),
    .rst(rst)
  );


endmodule
