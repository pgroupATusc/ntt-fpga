// NTT Accelerator

module NTT_Top #(
    parameter DATA_WIDTH_PER_INPUT = 28,
    parameter INPUT_PER_CYCLE = 64
  ) (
    inData,
    outData,
    in_start,
    out_start,
    clk,
    rst,
  );

  input clk, rst;

  input in_start[9:0];
  output logic out_start[9:0];

  input        [DATA_WIDTH_PER_INPUT-1:0] inData[INPUT_PER_CYCLE-1:0];
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_0_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_0_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_1_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_1_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_2_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_2_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_3_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_3_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_4_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_4_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_5_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_5_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_6_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_6_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_7_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_7_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_8_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_8_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_9_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_9_per_out[INPUT_PER_CYCLE-1:0];

  parameter [7:0] START_CYCLE[11] = {0, 7, 14, 21, 28, 35, 58, 82, 108, 138, 176};

  // TODO(Tian): stage 0 32 butterfly units
  butterfly #(
    .start(START_CYCLE[0]),
    .factors({66687, 58085086, 153619107, 41046131, 189026714, 70631961, 197498270, 125081754,
              54194127, 186938437, 218565763, 176985668, 66993197, 149817301, 44349942, 106663692,
              209875154, 265093046, 243595082, 40001367, 188637512, 130849588, 80900544, 41376169,
              74661667, 9521161, 117448591, 216779302, 67400723, 241368847, 190155959, 121954140}))
  stage_0_butterfly_0 (
    .x_in(inData[0]),
    .y_in(inData[1]),
    .x_out(stage_0_per_in[0]),
    .y_out(stage_0_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({69710552, 157049837, 29541109, 109238580, 176646986, 66294444, 4184358, 261365258,
              216344829, 157159811, 218464636, 109752985, 107013281, 83173794, 82066131, 127177690,
              211324969, 73580010, 262853884, 104968162, 241404981, 127320617, 96861137, 111883252,
              163120146, 164222678, 180135303, 222243486, 47960804, 11479903, 185458452, 14425613}))
  stage_0_butterfly_1 (
    .x_in(inData[2]),
    .y_in(inData[3]),
    .x_out(stage_0_per_in[2]),
    .y_out(stage_0_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({262755833, 25367770, 72606471, 131386739, 24152300, 113066699, 230614882, 212990958,
              83248807, 224274217, 56718282, 64307891, 80152118, 6554463, 249749550, 177333030,
              112928859, 103520242, 11377467, 212660495, 9977836, 248813222, 256522921, 42903438,
              243952581, 81165688, 13005428, 122372515, 127264350, 194452250, 97371131, 250007587}))
  stage_0_butterfly_2 (
    .x_in(inData[4]),
    .y_in(inData[5]),
    .x_out(stage_0_per_in[4]),
    .y_out(stage_0_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({256317058, 176574100, 196552678, 4087463, 197359850, 144888817, 116252651, 251186267,
              227177249, 37869546, 254559948, 80396852, 267404879, 243900215, 230038199, 186920055,
              183986337, 143442800, 77239454, 9418848, 136554761, 30998042, 234127283, 28513237,
              7407334, 185511309, 246139244, 207114911, 48499686, 132216843, 65241583, 13394971}))
  stage_0_butterfly_3 (
    .x_in(inData[6]),
    .y_in(inData[7]),
    .x_out(stage_0_per_in[6]),
    .y_out(stage_0_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({36785021, 116176624, 241027889, 2568552, 135965343, 220939348, 67459976, 156421542,
              53251080, 139206238, 37830528, 85925921, 250343614, 64508043, 92664685, 16229147,
              259190760, 5284602, 178626802, 34279912, 186026798, 229577517, 159848863, 132170867,
              118263349, 183471966, 188624074, 35688570, 133533317, 204610446, 96783518, 129161289}))
  stage_0_butterfly_4 (
    .x_in(inData[8]),
    .y_in(inData[9]),
    .x_out(stage_0_per_in[8]),
    .y_out(stage_0_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({70884448, 20380320, 62553766, 246330337, 17337072, 259358426, 221333762, 79007221,
              125436993, 165481068, 34758721, 76840577, 119165597, 143713813, 57880935, 159288788,
              185327331, 121708429, 26950622, 31628247, 116219557, 64402402, 86425411, 210629837,
              264754058, 160223263, 189299702, 38129962, 112174110, 148301509, 75689991, 181758089}))
  stage_0_butterfly_5 (
    .x_in(inData[10]),
    .y_in(inData[11]),
    .x_out(stage_0_per_in[10]),
    .y_out(stage_0_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({144486207, 33861678, 62424622, 171258656, 30978406, 191233099, 108814743, 200295213,
              240329350, 119553807, 17095567, 119820987, 125990181, 74620568, 195258296, 211474022,
              213018760, 217483488, 224076531, 124175107, 241147279, 43396787, 163686509, 267034870,
              21814275, 119858575, 233629950, 65363597, 61366355, 128923754, 207436891, 258398710}))
  stage_0_butterfly_6 (
    .x_in(inData[12]),
    .y_in(inData[13]),
    .x_out(stage_0_per_in[12]),
    .y_out(stage_0_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({4869479, 226423252, 240913336, 161193348, 7525756, 183816509, 45529198, 227631635,
              117082039, 85943438, 5742112, 55952036, 158362238, 114499544, 183015243, 224620084,
              98446051, 90415400, 202037642, 80852279, 219647998, 85610695, 35399020, 16387901,
              70993112, 56349189, 89363633, 72373951, 135336752, 211284483, 102019874, 212643172}))
  stage_0_butterfly_7 (
    .x_in(inData[14]),
    .y_in(inData[15]),
    .x_out(stage_0_per_in[14]),
    .y_out(stage_0_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({181036575, 15406607, 118216948, 28990836, 153827860, 152434516, 95356163, 190584784,
              104721465, 207179347, 195777196, 62694765, 192617727, 199997052, 185375251, 141917139,
              171269635, 66106013, 236173805, 48487396, 86222094, 64123411, 86412198, 29149935,
              67895486, 111028502, 220487343, 129596600, 126869459, 74346844, 115863951, 9083394}))
  stage_0_butterfly_8 (
    .x_in(inData[16]),
    .y_in(inData[17]),
    .x_out(stage_0_per_in[16]),
    .y_out(stage_0_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({164585197, 84197948, 162343477, 24580196, 112847505, 104494180, 239438610, 195751196,
              255042189, 27101256, 167135704, 178774268, 126420356, 60187882, 92935276, 201970932,
              242966976, 100723721, 113735821, 128081279, 209335538, 55000619, 40931981, 3906588,
              254651521, 6839312, 126673466, 35544064, 257856584, 240580313, 218254116, 28589493}))
  stage_0_butterfly_9 (
    .x_in(inData[18]),
    .y_in(inData[19]),
    .x_out(stage_0_per_in[18]),
    .y_out(stage_0_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({124689641, 12048336, 16967674, 165964934, 63479516, 264758616, 246348641, 12994463,
              151222684, 126817458, 15203085, 266062977, 158406994, 118812967, 231508432, 209775390,
              145325214, 115675578, 246040827, 131952477, 128639456, 174110644, 151896708, 248430418,
              43308742, 68558047, 186490797, 26451456, 227605745, 81924749, 100306740, 187430880}))
  stage_0_butterfly_10 (
    .x_in(inData[20]),
    .y_in(inData[21]),
    .x_out(stage_0_per_in[20]),
    .y_out(stage_0_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({236609676, 155632772, 208367077, 237702991, 192156570, 169217935, 111861272, 141932586,
              46680870, 4080689, 91771920, 64186729, 196972136, 24281843, 81641436, 120623833,
              224193580, 181657279, 114906207, 157158700, 66698835, 246446391, 15304900, 41918325,
              79432680, 35256934, 46133075, 228992312, 185850221, 34535827, 267892175, 94113816}))
  stage_0_butterfly_11 (
    .x_in(inData[22]),
    .y_in(inData[23]),
    .x_out(stage_0_per_in[22]),
    .y_out(stage_0_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({175181826, 25921170, 129053745, 59004276, 89839882, 119598304, 180106398, 75588758,
              94844905, 232035425, 76258087, 194631063, 129973973, 182519003, 13646129, 215427609,
              111161696, 182035415, 143397255, 175887545, 218411001, 242432529, 127510598, 210485515,
              214331009, 124878920, 181264550, 103427147, 239446376, 6261383, 100616259, 213513532}))
  stage_0_butterfly_12 (
    .x_in(inData[24]),
    .y_in(inData[25]),
    .x_out(stage_0_per_in[24]),
    .y_out(stage_0_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({53666796, 201841490, 250734390, 21867329, 195126393, 18807047, 154135831, 96098889,
              201750613, 56301526, 226796218, 75267274, 215876710, 86146205, 242906033, 106441080,
              51299486, 183906538, 186023395, 149121135, 37292607, 66456987, 127868408, 95362545,
              159083887, 124980045, 41512397, 216420108, 35769351, 177659362, 254862428, 175699854}))
  stage_0_butterfly_13 (
    .x_in(inData[26]),
    .y_in(inData[27]),
    .x_out(stage_0_per_in[26]),
    .y_out(stage_0_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({134572374, 54591848, 259641163, 266184237, 124903743, 243356346, 110349263, 217947353,
              260055946, 260941520, 39159482, 198451374, 188610091, 143647295, 16321430, 85861280,
              196727396, 4628244, 259902883, 176734838, 52172809, 88659311, 37689469, 246253529,
              263768524, 44002169, 153805373, 164064761, 16680201, 72006316, 104486975, 161494327}))
  stage_0_butterfly_14 (
    .x_in(inData[28]),
    .y_in(inData[29]),
    .x_out(stage_0_per_in[28]),
    .y_out(stage_0_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({251547338, 187954050, 9599856, 253615348, 145040924, 31515852, 75051406, 158367942,
              245518247, 147907047, 126638229, 197375798, 13677670, 208399648, 45577615, 102496219,
              259597052, 139662643, 140652682, 88068083, 22419281, 154457559, 209499403, 119681087,
              202709135, 11713205, 221869909, 187446019, 13905102, 61031492, 236043136, 81363847}))
  stage_0_butterfly_15 (
    .x_in(inData[30]),
    .y_in(inData[31]),
    .x_out(stage_0_per_in[30]),
    .y_out(stage_0_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({207692352, 171518128, 45213202, 231691713, 184120139, 79909455, 20654843, 22483780,
              241662912, 53018448, 29126603, 166849602, 242981970, 134488788, 215932651, 230537579,
              123744505, 13110486, 204305824, 124635721, 213462715, 188476710, 13136617, 134518349,
              22903087, 79252444, 34884345, 94872102, 110850189, 200589425, 7804022, 138643341}))
  stage_0_butterfly_16 (
    .x_in(inData[32]),
    .y_in(inData[33]),
    .x_out(stage_0_per_in[32]),
    .y_out(stage_0_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({255875272, 60493834, 199654780, 264692686, 222469354, 156023579, 164354184, 264722248,
              224632066, 42984958, 10057303, 19948338, 224618046, 78067214, 174707320, 111544693,
              42559975, 58402192, 135644103, 29014999, 248367053, 153843002, 52859373, 212200386,
              114169496, 261854403, 98181554, 251666562, 29380441, 205236983, 2705617, 214088558}))
  stage_0_butterfly_17 (
    .x_in(inData[34]),
    .y_in(inData[35]),
    .x_out(stage_0_per_in[34]),
    .y_out(stage_0_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({154212375, 14131216, 254000355, 248921617, 43817935, 181198907, 168908433, 9304145,
              255369977, 53103748, 127930513, 267667077, 18101390, 152808181, 144813234, 120419308,
              142863934, 121172029, 125480758, 205274966, 177181340, 1429580, 153907308, 198035948,
              124518160, 258225039, 107122996, 78535147, 90748831, 48447796, 210266721, 25148713}))
  stage_0_butterfly_18 (
    .x_in(inData[36]),
    .y_in(inData[37]),
    .x_out(stage_0_per_in[36]),
    .y_out(stage_0_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({5651134, 235215540, 65092548, 246972075, 205553550, 254205318, 219432305, 209423491,
              52761187, 77043356, 268253695, 243436973, 145663803, 207221115, 193252183, 178131021,
              153035867, 141410653, 209091203, 202016934, 105651679, 219873665, 130965208, 263341785,
              46629005, 119697484, 219164507, 200991325, 99140149, 169530517, 37489037, 233412603}))
  stage_0_butterfly_19 (
    .x_in(inData[38]),
    .y_in(inData[39]),
    .x_out(stage_0_per_in[38]),
    .y_out(stage_0_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({96644160, 238066757, 95745785, 94477870, 173093264, 20028125, 24122396, 145706676,
              130184658, 182490652, 176845896, 200245646, 75240990, 78372181, 175360485, 230913482,
              13214022, 72907110, 158913333, 144340508, 3731063, 193915015, 20163279, 143364478,
              124384681, 218119669, 8903594, 162610901, 224762304, 176649880, 101221270, 91136142}))
  stage_0_butterfly_20 (
    .x_in(inData[40]),
    .y_in(inData[41]),
    .x_out(stage_0_per_in[40]),
    .y_out(stage_0_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({208516738, 156384032, 38429557, 18485653, 107466416, 74839506, 76096071, 101664410,
              155494097, 83440545, 24169593, 214277734, 132749847, 15448747, 243480557, 232016200,
              200835165, 150529015, 218922070, 176876579, 241656403, 121678256, 199114532, 144387747,
              75455626, 237212534, 56848151, 189248627, 92098334, 234435452, 238700391, 35697312}))
  stage_0_butterfly_21 (
    .x_in(inData[42]),
    .y_in(inData[43]),
    .x_out(stage_0_per_in[42]),
    .y_out(stage_0_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({141475285, 122417419, 114175494, 187658742, 41031357, 82105625, 76495986, 78726832,
              204045920, 41015351, 184775632, 215044990, 216035935, 100034642, 187345691, 123869779,
              182322028, 172927150, 172413463, 226568978, 81774581, 126650083, 64059298, 200458300,
              229077055, 267701123, 116261862, 50041017, 114456140, 28569588, 12549924, 113970703}))
  stage_0_butterfly_22 (
    .x_in(inData[44]),
    .y_in(inData[45]),
    .x_out(stage_0_per_in[44]),
    .y_out(stage_0_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({250979164, 101235253, 219155874, 75430495, 127603059, 7373784, 150750886, 106279827,
              8437385, 241484731, 210367757, 50956256, 184194991, 88850354, 73886338, 202657965,
              222855093, 20476611, 117740425, 210930243, 159837268, 250769297, 1381761, 104273059,
              56672741, 15252454, 230462114, 260125445, 196403691, 179888950, 161018204, 228180092}))
  stage_0_butterfly_23 (
    .x_in(inData[46]),
    .y_in(inData[47]),
    .x_out(stage_0_per_in[46]),
    .y_out(stage_0_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({149046252, 249303130, 197016099, 127667482, 219408463, 90833651, 88694916, 154780521,
              152028008, 210835738, 91129770, 54694187, 233855133, 159375180, 89556414, 153057061,
              172630653, 229787934, 64197737, 174554842, 236960516, 144089543, 194834330, 182882105,
              50484120, 143928593, 77305748, 221852517, 60951044, 232958416, 185120175, 218263368}))
  stage_0_butterfly_24 (
    .x_in(inData[48]),
    .y_in(inData[49]),
    .x_out(stage_0_per_in[48]),
    .y_out(stage_0_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({82259521, 196076822, 208392312, 205950205, 194382796, 58882681, 226909804, 57420105,
              104225870, 265484036, 162889363, 101451720, 222836343, 146642358, 100770703, 94729012,
              253791818, 11727916, 114289273, 122009767, 206932975, 218155940, 246263559, 207289252,
              50021352, 22696094, 74643322, 33986901, 247062782, 3059556, 127281316, 202839194}))
  stage_0_butterfly_25 (
    .x_in(inData[50]),
    .y_in(inData[51]),
    .x_out(stage_0_per_in[50]),
    .y_out(stage_0_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({89494679, 172777377, 75161941, 173116375, 209076586, 33161823, 52952054, 79746145,
              219476260, 188253439, 217984510, 49412866, 263485445, 263389379, 184266218, 116815899,
              124256170, 236561162, 119485143, 59945410, 214979600, 214652925, 218479673, 242718809,
              125264465, 111988251, 77506253, 197145719, 122774092, 130025327, 220111512, 80477336}))
  stage_0_butterfly_26 (
    .x_in(inData[52]),
    .y_in(inData[53]),
    .x_out(stage_0_per_in[52]),
    .y_out(stage_0_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({108936038, 11247416, 12030631, 148728622, 139714595, 242696977, 232215778, 176645554,
              134032627, 253775510, 5933624, 204816575, 60114085, 101380813, 131659808, 40136402,
              41504705, 14923017, 1996702, 72665107, 203299319, 140980229, 185097589, 63912782,
              54250256, 172134458, 70728737, 37207751, 95857789, 202868018, 44186331, 172355039}))
  stage_0_butterfly_27 (
    .x_in(inData[54]),
    .y_in(inData[55]),
    .x_out(stage_0_per_in[54]),
    .y_out(stage_0_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({9453674, 122635188, 71023991, 7487276, 234963902, 99687432, 7289546, 195650024,
              232700332, 73305984, 76831465, 122925753, 136763023, 45684920, 170218646, 19111856,
              184394225, 34093582, 189966412, 6456449, 25932042, 207587513, 177566022, 148535761,
              114664154, 207578860, 69161829, 157107117, 14128368, 63900610, 126629575, 248049881}))
  stage_0_butterfly_28 (
    .x_in(inData[56]),
    .y_in(inData[57]),
    .x_out(stage_0_per_in[56]),
    .y_out(stage_0_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({149565630, 229646063, 32353046, 94417879, 223749061, 151510274, 175735543, 19569387,
              179997990, 268223107, 176150397, 146917464, 246670007, 220989018, 130341794, 245173438,
              168090046, 133543242, 36426289, 32769539, 33343400, 246049881, 190924029, 195750117,
              83665434, 79351768, 71466452, 132980811, 44753328, 15241225, 255807486, 100791881}))
  stage_0_butterfly_29 (
    .x_in(inData[58]),
    .y_in(inData[59]),
    .x_out(stage_0_per_in[58]),
    .y_out(stage_0_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({20490089, 172426762, 54291647, 83798709, 240846316, 252329804, 106939991, 39161232,
              62605527, 121709085, 194584338, 111058309, 189935724, 177655074, 239135625, 121236629,
              197999089, 85557225, 127312784, 233358957, 222818810, 65939487, 35608242, 217412044,
              66352780, 50385541, 203207502, 38583127, 178750844, 178548754, 259334239, 85449542}))
  stage_0_butterfly_30 (
    .x_in(inData[60]),
    .y_in(inData[61]),
    .x_out(stage_0_per_in[60]),
    .y_out(stage_0_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({198469359, 200880844, 107222748, 106713399, 94741987, 89730483, 92263376, 6208689,
              243959994, 132063071, 70296940, 91839141, 97932506, 117068649, 144316291, 258128862,
              244981517, 254780782, 75414331, 209997049, 103192680, 213843220, 241593066, 90431622,
              230254857, 92468150, 263850390, 231864746, 14195884, 180859208, 5071752, 86422302}))
  stage_0_butterfly_31 (
    .x_in(inData[62]),
    .y_in(inData[63]),
    .x_out(stage_0_per_in[62]),
    .y_out(stage_0_per_in[63]),
    .clk(clk),
    .rst(rst)
  );



  // TODO(Yang): stage 0 -> stage 1 permutation
  // FIXME: ignore butterfly units for now.
  stage_0_permutation #(
    .DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    .INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_0_1_per (
    .inData_0(stage_0_per_in[0]),
    .inData_1(stage_0_per_in[1]),
    .inData_2(stage_0_per_in[2]),
    .inData_3(stage_0_per_in[3]),
    .inData_4(stage_0_per_in[4]),
    .inData_5(stage_0_per_in[5]),
    .inData_6(stage_0_per_in[6]),
    .inData_7(stage_0_per_in[7]),
    .inData_8(stage_0_per_in[8]),
    .inData_9(stage_0_per_in[9]),
    .inData_10(stage_0_per_in[10]),
    .inData_11(stage_0_per_in[11]),
    .inData_12(stage_0_per_in[12]),
    .inData_13(stage_0_per_in[13]),
    .inData_14(stage_0_per_in[14]),
    .inData_15(stage_0_per_in[15]),
    .inData_16(stage_0_per_in[16]),
    .inData_17(stage_0_per_in[17]),
    .inData_18(stage_0_per_in[18]),
    .inData_19(stage_0_per_in[19]),
    .inData_20(stage_0_per_in[20]),
    .inData_21(stage_0_per_in[21]),
    .inData_22(stage_0_per_in[22]),
    .inData_23(stage_0_per_in[23]),
    .inData_24(stage_0_per_in[24]),
    .inData_25(stage_0_per_in[25]),
    .inData_26(stage_0_per_in[26]),
    .inData_27(stage_0_per_in[27]),
    .inData_28(stage_0_per_in[28]),
    .inData_29(stage_0_per_in[29]),
    .inData_30(stage_0_per_in[30]),
    .inData_31(stage_0_per_in[31]),
    .inData_32(stage_0_per_in[32]),
    .inData_33(stage_0_per_in[33]),
    .inData_34(stage_0_per_in[34]),
    .inData_35(stage_0_per_in[35]),
    .inData_36(stage_0_per_in[36]),
    .inData_37(stage_0_per_in[37]),
    .inData_38(stage_0_per_in[38]),
    .inData_39(stage_0_per_in[39]),
    .inData_40(stage_0_per_in[40]),
    .inData_41(stage_0_per_in[41]),
    .inData_42(stage_0_per_in[42]),
    .inData_43(stage_0_per_in[43]),
    .inData_44(stage_0_per_in[44]),
    .inData_45(stage_0_per_in[45]),
    .inData_46(stage_0_per_in[46]),
    .inData_47(stage_0_per_in[47]),
    .inData_48(stage_0_per_in[48]),
    .inData_49(stage_0_per_in[49]),
    .inData_50(stage_0_per_in[50]),
    .inData_51(stage_0_per_in[51]),
    .inData_52(stage_0_per_in[52]),
    .inData_53(stage_0_per_in[53]),
    .inData_54(stage_0_per_in[54]),
    .inData_55(stage_0_per_in[55]),
    .inData_56(stage_0_per_in[56]),
    .inData_57(stage_0_per_in[57]),
    .inData_58(stage_0_per_in[58]),
    .inData_59(stage_0_per_in[59]),
    .inData_60(stage_0_per_in[60]),
    .inData_61(stage_0_per_in[61]),
    .inData_62(stage_0_per_in[62]),
    .inData_63(stage_0_per_in[63]),
    .outData_0(stage_0_per_out[0]),
    .outData_1(stage_0_per_out[1]),
    .outData_2(stage_0_per_out[2]),
    .outData_3(stage_0_per_out[3]),
    .outData_4(stage_0_per_out[4]),
    .outData_5(stage_0_per_out[5]),
    .outData_6(stage_0_per_out[6]),
    .outData_7(stage_0_per_out[7]),
    .outData_8(stage_0_per_out[8]),
    .outData_9(stage_0_per_out[9]),
    .outData_10(stage_0_per_out[10]),
    .outData_11(stage_0_per_out[11]),
    .outData_12(stage_0_per_out[12]),
    .outData_13(stage_0_per_out[13]),
    .outData_14(stage_0_per_out[14]),
    .outData_15(stage_0_per_out[15]),
    .outData_16(stage_0_per_out[16]),
    .outData_17(stage_0_per_out[17]),
    .outData_18(stage_0_per_out[18]),
    .outData_19(stage_0_per_out[19]),
    .outData_20(stage_0_per_out[20]),
    .outData_21(stage_0_per_out[21]),
    .outData_22(stage_0_per_out[22]),
    .outData_23(stage_0_per_out[23]),
    .outData_24(stage_0_per_out[24]),
    .outData_25(stage_0_per_out[25]),
    .outData_26(stage_0_per_out[26]),
    .outData_27(stage_0_per_out[27]),
    .outData_28(stage_0_per_out[28]),
    .outData_29(stage_0_per_out[29]),
    .outData_30(stage_0_per_out[30]),
    .outData_31(stage_0_per_out[31]),
    .outData_32(stage_0_per_out[32]),
    .outData_33(stage_0_per_out[33]),
    .outData_34(stage_0_per_out[34]),
    .outData_35(stage_0_per_out[35]),
    .outData_36(stage_0_per_out[36]),
    .outData_37(stage_0_per_out[37]),
    .outData_38(stage_0_per_out[38]),
    .outData_39(stage_0_per_out[39]),
    .outData_40(stage_0_per_out[40]),
    .outData_41(stage_0_per_out[41]),
    .outData_42(stage_0_per_out[42]),
    .outData_43(stage_0_per_out[43]),
    .outData_44(stage_0_per_out[44]),
    .outData_45(stage_0_per_out[45]),
    .outData_46(stage_0_per_out[46]),
    .outData_47(stage_0_per_out[47]),
    .outData_48(stage_0_per_out[48]),
    .outData_49(stage_0_per_out[49]),
    .outData_50(stage_0_per_out[50]),
    .outData_51(stage_0_per_out[51]),
    .outData_52(stage_0_per_out[52]),
    .outData_53(stage_0_per_out[53]),
    .outData_54(stage_0_per_out[54]),
    .outData_55(stage_0_per_out[55]),
    .outData_56(stage_0_per_out[56]),
    .outData_57(stage_0_per_out[57]),
    .outData_58(stage_0_per_out[58]),
    .outData_59(stage_0_per_out[59]),
    .outData_60(stage_0_per_out[60]),
    .outData_61(stage_0_per_out[61]),
    .outData_62(stage_0_per_out[62]),
    .outData_63(stage_0_per_out[63]),
    .in_start(in_start[0]),
    .out_start(out_start[0]),
    .clk(clk),
    .rst(rst)
  );

  // TODO(Tian): stage 1 32 butterfly units
  butterfly #(
    .start(START_CYCLE[1]),
    .factors({153237233, 76624935, 137060289, 103368916, 180764097, 265109260, 138513718, 232173019,
              20917227, 227453822, 73099736, 168674209, 44888494, 135080569, 121414397, 261458154,
              174391063, 160856494, 43977927, 135902522, 56257750, 172655984, 2486257, 82483914,
              21253452, 99543252, 259302720, 267785378, 128052734, 244216061, 205242220, 20236367}))
  stage_1_butterfly_0 (
    .x_in(stage_0_per_out[0]),
    .y_in(stage_0_per_out[1]),
    .x_out(stage_1_per_in[0]),
    .y_out(stage_1_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({153237233, 76624935, 137060289, 103368916, 180764097, 265109260, 138513718, 232173019,
              20917227, 227453822, 73099736, 168674209, 44888494, 135080569, 121414397, 261458154,
              174391063, 160856494, 43977927, 135902522, 56257750, 172655984, 2486257, 82483914,
              21253452, 99543252, 259302720, 267785378, 128052734, 244216061, 205242220, 20236367}))
  stage_1_butterfly_1 (
    .x_in(stage_0_per_out[2]),
    .y_in(stage_0_per_out[3]),
    .x_out(stage_1_per_in[2]),
    .y_out(stage_1_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({83809662, 57946842, 46312994, 15655486, 172715743, 9793208, 160048836, 66337349,
              228243008, 56207397, 119878395, 42575603, 205934027, 59894768, 112070980, 159148996,
              89028484, 166334964, 134161265, 78767945, 21649526, 34932582, 112825183, 253487730,
              170100736, 36492987, 209643171, 228572460, 144648965, 232038388, 72369588, 171841734}))
  stage_1_butterfly_2 (
    .x_in(stage_0_per_out[4]),
    .y_in(stage_0_per_out[5]),
    .x_out(stage_1_per_in[4]),
    .y_out(stage_1_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({83809662, 57946842, 46312994, 15655486, 172715743, 9793208, 160048836, 66337349,
              228243008, 56207397, 119878395, 42575603, 205934027, 59894768, 112070980, 159148996,
              89028484, 166334964, 134161265, 78767945, 21649526, 34932582, 112825183, 253487730,
              170100736, 36492987, 209643171, 228572460, 144648965, 232038388, 72369588, 171841734}))
  stage_1_butterfly_3 (
    .x_in(stage_0_per_out[6]),
    .y_in(stage_0_per_out[7]),
    .x_out(stage_1_per_in[6]),
    .y_out(stage_1_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({257723260, 25278905, 164865927, 121608761, 245986816, 85740049, 46282885, 82779345,
              156534179, 74931497, 226025718, 255818084, 76313029, 242717180, 249947221, 262630184,
              113006603, 175949223, 187381670, 188535281, 234775081, 90701762, 217359458, 94178347,
              248946430, 267860193, 191242693, 44896056, 10943590, 136898494, 87202745, 237616434}))
  stage_1_butterfly_4 (
    .x_in(stage_0_per_out[8]),
    .y_in(stage_0_per_out[9]),
    .x_out(stage_1_per_in[8]),
    .y_out(stage_1_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({257723260, 25278905, 164865927, 121608761, 245986816, 85740049, 46282885, 82779345,
              156534179, 74931497, 226025718, 255818084, 76313029, 242717180, 249947221, 262630184,
              113006603, 175949223, 187381670, 188535281, 234775081, 90701762, 217359458, 94178347,
              248946430, 267860193, 191242693, 44896056, 10943590, 136898494, 87202745, 237616434}))
  stage_1_butterfly_5 (
    .x_in(stage_0_per_out[10]),
    .y_in(stage_0_per_out[11]),
    .x_out(stage_1_per_in[10]),
    .y_out(stage_1_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({267008435, 65803974, 198352904, 133573372, 53126225, 211646222, 185175266, 233083676,
              207021189, 219133933, 78273516, 67241659, 138629310, 143811089, 13228372, 122025398,
              18793692, 155613159, 45457492, 116513948, 99899421, 31964447, 198957507, 116527240,
              53025186, 232740066, 146205579, 50523873, 264322432, 16351380, 159987098, 165584204}))
  stage_1_butterfly_6 (
    .x_in(stage_0_per_out[12]),
    .y_in(stage_0_per_out[13]),
    .x_out(stage_1_per_in[12]),
    .y_out(stage_1_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({267008435, 65803974, 198352904, 133573372, 53126225, 211646222, 185175266, 233083676,
              207021189, 219133933, 78273516, 67241659, 138629310, 143811089, 13228372, 122025398,
              18793692, 155613159, 45457492, 116513948, 99899421, 31964447, 198957507, 116527240,
              53025186, 232740066, 146205579, 50523873, 264322432, 16351380, 159987098, 165584204}))
  stage_1_butterfly_7 (
    .x_in(stage_0_per_out[14]),
    .y_in(stage_0_per_out[15]),
    .x_out(stage_1_per_in[14]),
    .y_out(stage_1_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({181617487, 5445105, 167645260, 266777383, 215525211, 210373784, 69017626, 193451294,
              243047656, 211824237, 5267255, 206844979, 18433789, 40915578, 12912005, 139742686,
              83977288, 125713617, 62456195, 251672258, 127163336, 74458128, 175710456, 230865684,
              176911171, 151857114, 146399832, 169792793, 44047649, 45355620, 205604517, 129677075}))
  stage_1_butterfly_8 (
    .x_in(stage_0_per_out[16]),
    .y_in(stage_0_per_out[17]),
    .x_out(stage_1_per_in[16]),
    .y_out(stage_1_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({181617487, 5445105, 167645260, 266777383, 215525211, 210373784, 69017626, 193451294,
              243047656, 211824237, 5267255, 206844979, 18433789, 40915578, 12912005, 139742686,
              83977288, 125713617, 62456195, 251672258, 127163336, 74458128, 175710456, 230865684,
              176911171, 151857114, 146399832, 169792793, 44047649, 45355620, 205604517, 129677075}))
  stage_1_butterfly_9 (
    .x_in(stage_0_per_out[18]),
    .y_in(stage_0_per_out[19]),
    .x_out(stage_1_per_in[18]),
    .y_out(stage_1_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({3395282, 36620312, 77119896, 195181845, 249311139, 87492030, 108319109, 129694458,
              19700796, 62513408, 199055975, 215085706, 7301415, 11850588, 116257755, 133565368,
              194684542, 157839041, 64830196, 17682401, 43819650, 236272786, 12286825, 182803613,
              94436408, 238832783, 84798700, 226834391, 209708523, 70944317, 141562255, 133273987}))
  stage_1_butterfly_10 (
    .x_in(stage_0_per_out[20]),
    .y_in(stage_0_per_out[21]),
    .x_out(stage_1_per_in[20]),
    .y_out(stage_1_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({3395282, 36620312, 77119896, 195181845, 249311139, 87492030, 108319109, 129694458,
              19700796, 62513408, 199055975, 215085706, 7301415, 11850588, 116257755, 133565368,
              194684542, 157839041, 64830196, 17682401, 43819650, 236272786, 12286825, 182803613,
              94436408, 238832783, 84798700, 226834391, 209708523, 70944317, 141562255, 133273987}))
  stage_1_butterfly_11 (
    .x_in(stage_0_per_out[22]),
    .y_in(stage_0_per_out[23]),
    .x_out(stage_1_per_in[22]),
    .y_out(stage_1_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({66412546, 17758040, 69205492, 105793954, 224922683, 98139687, 244004517, 40741603,
              213678985, 226759664, 91397014, 94686133, 74472522, 112360014, 47531240, 203850982,
              60051251, 50162577, 219484262, 232847226, 16652121, 196018390, 56132215, 90149574,
              50083600, 154298223, 106743034, 139044757, 149788353, 97163404, 265496406, 77783793}))
  stage_1_butterfly_12 (
    .x_in(stage_0_per_out[24]),
    .y_in(stage_0_per_out[25]),
    .x_out(stage_1_per_in[24]),
    .y_out(stage_1_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({66412546, 17758040, 69205492, 105793954, 224922683, 98139687, 244004517, 40741603,
              213678985, 226759664, 91397014, 94686133, 74472522, 112360014, 47531240, 203850982,
              60051251, 50162577, 219484262, 232847226, 16652121, 196018390, 56132215, 90149574,
              50083600, 154298223, 106743034, 139044757, 149788353, 97163404, 265496406, 77783793}))
  stage_1_butterfly_13 (
    .x_in(stage_0_per_out[26]),
    .y_in(stage_0_per_out[27]),
    .x_out(stage_1_per_in[26]),
    .y_out(stage_1_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({3341663, 157386503, 190540901, 229954056, 90687088, 226981541, 211982342, 175990762,
              18338102, 260110386, 107024087, 81838336, 136710753, 255463943, 263001722, 101579460,
              163823140, 160539079, 2017030, 86776671, 228715598, 25360705, 126413069, 19904170,
              77804235, 120080647, 238468357, 92441360, 78612624, 254842567, 172401093, 79230237}))
  stage_1_butterfly_14 (
    .x_in(stage_0_per_out[28]),
    .y_in(stage_0_per_out[29]),
    .x_out(stage_1_per_in[28]),
    .y_out(stage_1_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({3341663, 157386503, 190540901, 229954056, 90687088, 226981541, 211982342, 175990762,
              18338102, 260110386, 107024087, 81838336, 136710753, 255463943, 263001722, 101579460,
              163823140, 160539079, 2017030, 86776671, 228715598, 25360705, 126413069, 19904170,
              77804235, 120080647, 238468357, 92441360, 78612624, 254842567, 172401093, 79230237}))
  stage_1_butterfly_15 (
    .x_in(stage_0_per_out[30]),
    .y_in(stage_0_per_out[31]),
    .x_out(stage_1_per_in[30]),
    .y_out(stage_1_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({165180840, 99012968, 100343421, 29594281, 167181901, 94741537, 243339369, 262368251,
              146639516, 164079161, 84700854, 46197346, 259533807, 193174373, 64771890, 73072346,
              38252193, 81263879, 217210388, 102698816, 133952844, 202480866, 259164217, 244022079,
              108831626, 121145061, 23442787, 267017218, 195692414, 212728405, 231354349, 3021514}))
  stage_1_butterfly_16 (
    .x_in(stage_0_per_out[32]),
    .y_in(stage_0_per_out[33]),
    .x_out(stage_1_per_in[32]),
    .y_out(stage_1_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({165180840, 99012968, 100343421, 29594281, 167181901, 94741537, 243339369, 262368251,
              146639516, 164079161, 84700854, 46197346, 259533807, 193174373, 64771890, 73072346,
              38252193, 81263879, 217210388, 102698816, 133952844, 202480866, 259164217, 244022079,
              108831626, 121145061, 23442787, 267017218, 195692414, 212728405, 231354349, 3021514}))
  stage_1_butterfly_17 (
    .x_in(stage_0_per_out[34]),
    .y_in(stage_0_per_out[35]),
    .x_out(stage_1_per_in[34]),
    .y_out(stage_1_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({168373202, 159491687, 73071114, 255737752, 156837559, 58491201, 244423105, 102243739,
              100611174, 1592710, 178382895, 189033696, 237395333, 164473684, 10310370, 72509307,
              54714468, 266378632, 98410858, 238590283, 107503597, 62027985, 122609533, 173513151,
              21582278, 107940029, 8748458, 7376627, 108164959, 113049121, 154317057, 34052825}))
  stage_1_butterfly_18 (
    .x_in(stage_0_per_out[36]),
    .y_in(stage_0_per_out[37]),
    .x_out(stage_1_per_in[36]),
    .y_out(stage_1_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({168373202, 159491687, 73071114, 255737752, 156837559, 58491201, 244423105, 102243739,
              100611174, 1592710, 178382895, 189033696, 237395333, 164473684, 10310370, 72509307,
              54714468, 266378632, 98410858, 238590283, 107503597, 62027985, 122609533, 173513151,
              21582278, 107940029, 8748458, 7376627, 108164959, 113049121, 154317057, 34052825}))
  stage_1_butterfly_19 (
    .x_in(stage_0_per_out[38]),
    .y_in(stage_0_per_out[39]),
    .x_out(stage_1_per_in[38]),
    .y_out(stage_1_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({4457103, 121355275, 236209279, 79121706, 75689102, 247714871, 128011618, 142807968,
              259719559, 67784869, 169092523, 94341361, 255478273, 2204580, 263649093, 12817079,
              50606491, 122969043, 202871094, 248922055, 214937778, 207877484, 201160126, 149904904,
              110378476, 70033082, 195152646, 104557844, 86359417, 39337018, 240930884, 128159746}))
  stage_1_butterfly_20 (
    .x_in(stage_0_per_out[40]),
    .y_in(stage_0_per_out[41]),
    .x_out(stage_1_per_in[40]),
    .y_out(stage_1_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({4457103, 121355275, 236209279, 79121706, 75689102, 247714871, 128011618, 142807968,
              259719559, 67784869, 169092523, 94341361, 255478273, 2204580, 263649093, 12817079,
              50606491, 122969043, 202871094, 248922055, 214937778, 207877484, 201160126, 149904904,
              110378476, 70033082, 195152646, 104557844, 86359417, 39337018, 240930884, 128159746}))
  stage_1_butterfly_21 (
    .x_in(stage_0_per_out[42]),
    .y_in(stage_0_per_out[43]),
    .x_out(stage_1_per_in[42]),
    .y_out(stage_1_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({248328138, 112174557, 12711531, 230871518, 254234203, 128995628, 161607031, 118444917,
              218195682, 148649408, 217993137, 148479452, 82321748, 24036023, 187988754, 132747224,
              184464011, 173577844, 1807449, 120217110, 86350556, 118320134, 188526794, 184177651,
              115050087, 186476418, 207530748, 7226699, 1855205, 7280660, 189909138, 123018041}))
  stage_1_butterfly_22 (
    .x_in(stage_0_per_out[44]),
    .y_in(stage_0_per_out[45]),
    .x_out(stage_1_per_in[44]),
    .y_out(stage_1_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({248328138, 112174557, 12711531, 230871518, 254234203, 128995628, 161607031, 118444917,
              218195682, 148649408, 217993137, 148479452, 82321748, 24036023, 187988754, 132747224,
              184464011, 173577844, 1807449, 120217110, 86350556, 118320134, 188526794, 184177651,
              115050087, 186476418, 207530748, 7226699, 1855205, 7280660, 189909138, 123018041}))
  stage_1_butterfly_23 (
    .x_in(stage_0_per_out[46]),
    .y_in(stage_0_per_out[47]),
    .x_out(stage_1_per_in[46]),
    .y_out(stage_1_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({207769332, 36213609, 34402629, 136179523, 120466187, 184522009, 246741831, 135921552,
              62094530, 259895089, 234786570, 64464693, 127918992, 100027171, 263648524, 241071152,
              248251528, 133098101, 73481957, 198043993, 81414740, 209744644, 187208958, 190453366,
              30998914, 32319537, 263725948, 54916848, 245372433, 128297265, 110720332, 23586243}))
  stage_1_butterfly_24 (
    .x_in(stage_0_per_out[48]),
    .y_in(stage_0_per_out[49]),
    .x_out(stage_1_per_in[48]),
    .y_out(stage_1_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({207769332, 36213609, 34402629, 136179523, 120466187, 184522009, 246741831, 135921552,
              62094530, 259895089, 234786570, 64464693, 127918992, 100027171, 263648524, 241071152,
              248251528, 133098101, 73481957, 198043993, 81414740, 209744644, 187208958, 190453366,
              30998914, 32319537, 263725948, 54916848, 245372433, 128297265, 110720332, 23586243}))
  stage_1_butterfly_25 (
    .x_in(stage_0_per_out[50]),
    .y_in(stage_0_per_out[51]),
    .x_out(stage_1_per_in[50]),
    .y_out(stage_1_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({164728317, 115053845, 110055875, 145831337, 204707946, 101783683, 212788230, 218380292,
              209780385, 54393228, 92902456, 174856430, 19817676, 98445813, 141267184, 209154967,
              222249559, 144502563, 84669572, 139101859, 104121890, 121712648, 26068775, 104215821,
              2487567, 216819035, 105443909, 97171493, 134561032, 138215130, 120261431, 248732744}))
  stage_1_butterfly_26 (
    .x_in(stage_0_per_out[52]),
    .y_in(stage_0_per_out[53]),
    .x_out(stage_1_per_in[52]),
    .y_out(stage_1_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({164728317, 115053845, 110055875, 145831337, 204707946, 101783683, 212788230, 218380292,
              209780385, 54393228, 92902456, 174856430, 19817676, 98445813, 141267184, 209154967,
              222249559, 144502563, 84669572, 139101859, 104121890, 121712648, 26068775, 104215821,
              2487567, 216819035, 105443909, 97171493, 134561032, 138215130, 120261431, 248732744}))
  stage_1_butterfly_27 (
    .x_in(stage_0_per_out[54]),
    .y_in(stage_0_per_out[55]),
    .x_out(stage_1_per_in[54]),
    .y_out(stage_1_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({206116619, 151297332, 128589211, 45842328, 268043824, 236829199, 236528116, 17642100,
              58671364, 183613005, 107152911, 55222727, 158067861, 113269084, 145317914, 37377133,
              18205961, 212287973, 33096679, 102230592, 189044804, 23328014, 863665, 209112367,
              148051010, 256834872, 211201491, 93757293, 187172755, 159978713, 158914825, 263207998}))
  stage_1_butterfly_28 (
    .x_in(stage_0_per_out[56]),
    .y_in(stage_0_per_out[57]),
    .x_out(stage_1_per_in[56]),
    .y_out(stage_1_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({206116619, 151297332, 128589211, 45842328, 268043824, 236829199, 236528116, 17642100,
              58671364, 183613005, 107152911, 55222727, 158067861, 113269084, 145317914, 37377133,
              18205961, 212287973, 33096679, 102230592, 189044804, 23328014, 863665, 209112367,
              148051010, 256834872, 211201491, 93757293, 187172755, 159978713, 158914825, 263207998}))
  stage_1_butterfly_29 (
    .x_in(stage_0_per_out[58]),
    .y_in(stage_0_per_out[59]),
    .x_out(stage_1_per_in[58]),
    .y_out(stage_1_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({207047180, 126749676, 142941966, 187867192, 123335487, 183590673, 174290656, 31243956,
              23776027, 94206887, 92770973, 12591284, 122455193, 118946466, 189816962, 212425161,
              163197321, 107138937, 77536776, 62688241, 58903295, 6257752, 197065781, 6828726,
              201787732, 43000087, 10967191, 75993973, 145056180, 6760936, 51838504, 55947412}))
  stage_1_butterfly_30 (
    .x_in(stage_0_per_out[60]),
    .y_in(stage_0_per_out[61]),
    .x_out(stage_1_per_in[60]),
    .y_out(stage_1_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({207047180, 126749676, 142941966, 187867192, 123335487, 183590673, 174290656, 31243956,
              23776027, 94206887, 92770973, 12591284, 122455193, 118946466, 189816962, 212425161,
              163197321, 107138937, 77536776, 62688241, 58903295, 6257752, 197065781, 6828726,
              201787732, 43000087, 10967191, 75993973, 145056180, 6760936, 51838504, 55947412}))
  stage_1_butterfly_31 (
    .x_in(stage_0_per_out[62]),
    .y_in(stage_0_per_out[63]),
    .x_out(stage_1_per_in[62]),
    .y_out(stage_1_per_in[63]),
    .clk(clk),
    .rst(rst)
  );



  
  // TODO(Yang): stage 1 -> stage 2 permutation
  // FIXME: ignore butterfly units for now.
  stage_1_permutation #(
    .DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    .INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_1_2_per (
    .inData_0(stage_1_per_in[0]),
    .inData_1(stage_1_per_in[1]),
    .inData_2(stage_1_per_in[2]),
    .inData_3(stage_1_per_in[3]),
    .inData_4(stage_1_per_in[4]),
    .inData_5(stage_1_per_in[5]),
    .inData_6(stage_1_per_in[6]),
    .inData_7(stage_1_per_in[7]),
    .inData_8(stage_1_per_in[8]),
    .inData_9(stage_1_per_in[9]),
    .inData_10(stage_1_per_in[10]),
    .inData_11(stage_1_per_in[11]),
    .inData_12(stage_1_per_in[12]),
    .inData_13(stage_1_per_in[13]),
    .inData_14(stage_1_per_in[14]),
    .inData_15(stage_1_per_in[15]),
    .inData_16(stage_1_per_in[16]),
    .inData_17(stage_1_per_in[17]),
    .inData_18(stage_1_per_in[18]),
    .inData_19(stage_1_per_in[19]),
    .inData_20(stage_1_per_in[20]),
    .inData_21(stage_1_per_in[21]),
    .inData_22(stage_1_per_in[22]),
    .inData_23(stage_1_per_in[23]),
    .inData_24(stage_1_per_in[24]),
    .inData_25(stage_1_per_in[25]),
    .inData_26(stage_1_per_in[26]),
    .inData_27(stage_1_per_in[27]),
    .inData_28(stage_1_per_in[28]),
    .inData_29(stage_1_per_in[29]),
    .inData_30(stage_1_per_in[30]),
    .inData_31(stage_1_per_in[31]),
    .inData_32(stage_1_per_in[32]),
    .inData_33(stage_1_per_in[33]),
    .inData_34(stage_1_per_in[34]),
    .inData_35(stage_1_per_in[35]),
    .inData_36(stage_1_per_in[36]),
    .inData_37(stage_1_per_in[37]),
    .inData_38(stage_1_per_in[38]),
    .inData_39(stage_1_per_in[39]),
    .inData_40(stage_1_per_in[40]),
    .inData_41(stage_1_per_in[41]),
    .inData_42(stage_1_per_in[42]),
    .inData_43(stage_1_per_in[43]),
    .inData_44(stage_1_per_in[44]),
    .inData_45(stage_1_per_in[45]),
    .inData_46(stage_1_per_in[46]),
    .inData_47(stage_1_per_in[47]),
    .inData_48(stage_1_per_in[48]),
    .inData_49(stage_1_per_in[49]),
    .inData_50(stage_1_per_in[50]),
    .inData_51(stage_1_per_in[51]),
    .inData_52(stage_1_per_in[52]),
    .inData_53(stage_1_per_in[53]),
    .inData_54(stage_1_per_in[54]),
    .inData_55(stage_1_per_in[55]),
    .inData_56(stage_1_per_in[56]),
    .inData_57(stage_1_per_in[57]),
    .inData_58(stage_1_per_in[58]),
    .inData_59(stage_1_per_in[59]),
    .inData_60(stage_1_per_in[60]),
    .inData_61(stage_1_per_in[61]),
    .inData_62(stage_1_per_in[62]),
    .inData_63(stage_1_per_in[63]),
    .outData_0(stage_1_per_out[0]),
    .outData_1(stage_1_per_out[1]),
    .outData_2(stage_1_per_out[2]),
    .outData_3(stage_1_per_out[3]),
    .outData_4(stage_1_per_out[4]),
    .outData_5(stage_1_per_out[5]),
    .outData_6(stage_1_per_out[6]),
    .outData_7(stage_1_per_out[7]),
    .outData_8(stage_1_per_out[8]),
    .outData_9(stage_1_per_out[9]),
    .outData_10(stage_1_per_out[10]),
    .outData_11(stage_1_per_out[11]),
    .outData_12(stage_1_per_out[12]),
    .outData_13(stage_1_per_out[13]),
    .outData_14(stage_1_per_out[14]),
    .outData_15(stage_1_per_out[15]),
    .outData_16(stage_1_per_out[16]),
    .outData_17(stage_1_per_out[17]),
    .outData_18(stage_1_per_out[18]),
    .outData_19(stage_1_per_out[19]),
    .outData_20(stage_1_per_out[20]),
    .outData_21(stage_1_per_out[21]),
    .outData_22(stage_1_per_out[22]),
    .outData_23(stage_1_per_out[23]),
    .outData_24(stage_1_per_out[24]),
    .outData_25(stage_1_per_out[25]),
    .outData_26(stage_1_per_out[26]),
    .outData_27(stage_1_per_out[27]),
    .outData_28(stage_1_per_out[28]),
    .outData_29(stage_1_per_out[29]),
    .outData_30(stage_1_per_out[30]),
    .outData_31(stage_1_per_out[31]),
    .outData_32(stage_1_per_out[32]),
    .outData_33(stage_1_per_out[33]),
    .outData_34(stage_1_per_out[34]),
    .outData_35(stage_1_per_out[35]),
    .outData_36(stage_1_per_out[36]),
    .outData_37(stage_1_per_out[37]),
    .outData_38(stage_1_per_out[38]),
    .outData_39(stage_1_per_out[39]),
    .outData_40(stage_1_per_out[40]),
    .outData_41(stage_1_per_out[41]),
    .outData_42(stage_1_per_out[42]),
    .outData_43(stage_1_per_out[43]),
    .outData_44(stage_1_per_out[44]),
    .outData_45(stage_1_per_out[45]),
    .outData_46(stage_1_per_out[46]),
    .outData_47(stage_1_per_out[47]),
    .outData_48(stage_1_per_out[48]),
    .outData_49(stage_1_per_out[49]),
    .outData_50(stage_1_per_out[50]),
    .outData_51(stage_1_per_out[51]),
    .outData_52(stage_1_per_out[52]),
    .outData_53(stage_1_per_out[53]),
    .outData_54(stage_1_per_out[54]),
    .outData_55(stage_1_per_out[55]),
    .outData_56(stage_1_per_out[56]),
    .outData_57(stage_1_per_out[57]),
    .outData_58(stage_1_per_out[58]),
    .outData_59(stage_1_per_out[59]),
    .outData_60(stage_1_per_out[60]),
    .outData_61(stage_1_per_out[61]),
    .outData_62(stage_1_per_out[62]),
    .outData_63(stage_1_per_out[63]),
    .in_start(in_start[1]),
    .out_start(out_start[1]),
    .clk(clk),
    .rst(rst)
  );


  // TODO(Tian): stage 2 32 butterfly units
  butterfly #(
    .start(START_CYCLE[2]),
    .factors({184644727, 171051327, 43104106, 224225395, 196522490, 167366585, 218147185, 213835479,
              193915204, 165350229, 206705681, 117507527, 242516310, 158168844, 165872957, 261795000,
              98085790, 67225153, 42355602, 28242170, 186863562, 259958064, 109479656, 182702557,
              242425786, 131304314, 82155735, 55609416, 141424302, 118377542, 92160417, 56246211}))
  stage_2_butterfly_0 (
    .x_in(stage_1_per_out[0]),
    .y_in(stage_1_per_out[1]),
    .x_out(stage_2_per_in[0]),
    .y_out(stage_2_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({184644727, 171051327, 43104106, 224225395, 196522490, 167366585, 218147185, 213835479,
              193915204, 165350229, 206705681, 117507527, 242516310, 158168844, 165872957, 261795000,
              98085790, 67225153, 42355602, 28242170, 186863562, 259958064, 109479656, 182702557,
              242425786, 131304314, 82155735, 55609416, 141424302, 118377542, 92160417, 56246211}))
  stage_2_butterfly_1 (
    .x_in(stage_1_per_out[2]),
    .y_in(stage_1_per_out[3]),
    .x_out(stage_2_per_in[2]),
    .y_out(stage_2_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({184644727, 171051327, 43104106, 224225395, 196522490, 167366585, 218147185, 213835479,
              193915204, 165350229, 206705681, 117507527, 242516310, 158168844, 165872957, 261795000,
              98085790, 67225153, 42355602, 28242170, 186863562, 259958064, 109479656, 182702557,
              242425786, 131304314, 82155735, 55609416, 141424302, 118377542, 92160417, 56246211}))
  stage_2_butterfly_2 (
    .x_in(stage_1_per_out[4]),
    .y_in(stage_1_per_out[5]),
    .x_out(stage_2_per_in[4]),
    .y_out(stage_2_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({184644727, 171051327, 43104106, 224225395, 196522490, 167366585, 218147185, 213835479,
              193915204, 165350229, 206705681, 117507527, 242516310, 158168844, 165872957, 261795000,
              98085790, 67225153, 42355602, 28242170, 186863562, 259958064, 109479656, 182702557,
              242425786, 131304314, 82155735, 55609416, 141424302, 118377542, 92160417, 56246211}))
  stage_2_butterfly_3 (
    .x_in(stage_1_per_out[6]),
    .y_in(stage_1_per_out[7]),
    .x_out(stage_2_per_in[6]),
    .y_out(stage_2_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({255286072, 173118058, 185138250, 134269022, 222861227, 200399539, 82684352, 69584498,
              87202272, 29987725, 21739535, 171362072, 119169851, 215146927, 244477824, 26067051,
              135886841, 160841949, 135618975, 157966005, 210795202, 14568946, 82934386, 100123291,
              251384491, 40550456, 262464837, 217383280, 206252403, 199810586, 129576773, 32087335}))
  stage_2_butterfly_4 (
    .x_in(stage_1_per_out[8]),
    .y_in(stage_1_per_out[9]),
    .x_out(stage_2_per_in[8]),
    .y_out(stage_2_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({255286072, 173118058, 185138250, 134269022, 222861227, 200399539, 82684352, 69584498,
              87202272, 29987725, 21739535, 171362072, 119169851, 215146927, 244477824, 26067051,
              135886841, 160841949, 135618975, 157966005, 210795202, 14568946, 82934386, 100123291,
              251384491, 40550456, 262464837, 217383280, 206252403, 199810586, 129576773, 32087335}))
  stage_2_butterfly_5 (
    .x_in(stage_1_per_out[10]),
    .y_in(stage_1_per_out[11]),
    .x_out(stage_2_per_in[10]),
    .y_out(stage_2_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({255286072, 173118058, 185138250, 134269022, 222861227, 200399539, 82684352, 69584498,
              87202272, 29987725, 21739535, 171362072, 119169851, 215146927, 244477824, 26067051,
              135886841, 160841949, 135618975, 157966005, 210795202, 14568946, 82934386, 100123291,
              251384491, 40550456, 262464837, 217383280, 206252403, 199810586, 129576773, 32087335}))
  stage_2_butterfly_6 (
    .x_in(stage_1_per_out[12]),
    .y_in(stage_1_per_out[13]),
    .x_out(stage_2_per_in[12]),
    .y_out(stage_2_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({255286072, 173118058, 185138250, 134269022, 222861227, 200399539, 82684352, 69584498,
              87202272, 29987725, 21739535, 171362072, 119169851, 215146927, 244477824, 26067051,
              135886841, 160841949, 135618975, 157966005, 210795202, 14568946, 82934386, 100123291,
              251384491, 40550456, 262464837, 217383280, 206252403, 199810586, 129576773, 32087335}))
  stage_2_butterfly_7 (
    .x_in(stage_1_per_out[14]),
    .y_in(stage_1_per_out[15]),
    .x_out(stage_2_per_in[14]),
    .y_out(stage_2_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({158466952, 196328787, 34971158, 81527994, 174900371, 32260862, 249146534, 233514072,
              47375162, 124400051, 161171966, 202776751, 218694662, 201863951, 158727274, 209583375,
              102915173, 134877507, 169508713, 23405380, 100229847, 160254284, 63079505, 244763177,
              40158424, 181468172, 77389872, 219312182, 9842125, 67321994, 207821787, 262540431}))
  stage_2_butterfly_8 (
    .x_in(stage_1_per_out[16]),
    .y_in(stage_1_per_out[17]),
    .x_out(stage_2_per_in[16]),
    .y_out(stage_2_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({158466952, 196328787, 34971158, 81527994, 174900371, 32260862, 249146534, 233514072,
              47375162, 124400051, 161171966, 202776751, 218694662, 201863951, 158727274, 209583375,
              102915173, 134877507, 169508713, 23405380, 100229847, 160254284, 63079505, 244763177,
              40158424, 181468172, 77389872, 219312182, 9842125, 67321994, 207821787, 262540431}))
  stage_2_butterfly_9 (
    .x_in(stage_1_per_out[18]),
    .y_in(stage_1_per_out[19]),
    .x_out(stage_2_per_in[18]),
    .y_out(stage_2_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({158466952, 196328787, 34971158, 81527994, 174900371, 32260862, 249146534, 233514072,
              47375162, 124400051, 161171966, 202776751, 218694662, 201863951, 158727274, 209583375,
              102915173, 134877507, 169508713, 23405380, 100229847, 160254284, 63079505, 244763177,
              40158424, 181468172, 77389872, 219312182, 9842125, 67321994, 207821787, 262540431}))
  stage_2_butterfly_10 (
    .x_in(stage_1_per_out[20]),
    .y_in(stage_1_per_out[21]),
    .x_out(stage_2_per_in[20]),
    .y_out(stage_2_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({158466952, 196328787, 34971158, 81527994, 174900371, 32260862, 249146534, 233514072,
              47375162, 124400051, 161171966, 202776751, 218694662, 201863951, 158727274, 209583375,
              102915173, 134877507, 169508713, 23405380, 100229847, 160254284, 63079505, 244763177,
              40158424, 181468172, 77389872, 219312182, 9842125, 67321994, 207821787, 262540431}))
  stage_2_butterfly_11 (
    .x_in(stage_1_per_out[22]),
    .y_in(stage_1_per_out[23]),
    .x_out(stage_2_per_in[22]),
    .y_out(stage_2_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({160807241, 177340471, 199876762, 125267062, 260909397, 229100654, 1562592, 55567611,
              43575145, 252241817, 237438985, 42585458, 129101436, 60072008, 1613379, 130696933,
              99187435, 250508912, 77981460, 178386996, 181295312, 64884498, 56094099, 13458851,
              20857483, 27056737, 114486793, 196771169, 61345534, 66242139, 151095818, 168977833}))
  stage_2_butterfly_12 (
    .x_in(stage_1_per_out[24]),
    .y_in(stage_1_per_out[25]),
    .x_out(stage_2_per_in[24]),
    .y_out(stage_2_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({160807241, 177340471, 199876762, 125267062, 260909397, 229100654, 1562592, 55567611,
              43575145, 252241817, 237438985, 42585458, 129101436, 60072008, 1613379, 130696933,
              99187435, 250508912, 77981460, 178386996, 181295312, 64884498, 56094099, 13458851,
              20857483, 27056737, 114486793, 196771169, 61345534, 66242139, 151095818, 168977833}))
  stage_2_butterfly_13 (
    .x_in(stage_1_per_out[26]),
    .y_in(stage_1_per_out[27]),
    .x_out(stage_2_per_in[26]),
    .y_out(stage_2_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({160807241, 177340471, 199876762, 125267062, 260909397, 229100654, 1562592, 55567611,
              43575145, 252241817, 237438985, 42585458, 129101436, 60072008, 1613379, 130696933,
              99187435, 250508912, 77981460, 178386996, 181295312, 64884498, 56094099, 13458851,
              20857483, 27056737, 114486793, 196771169, 61345534, 66242139, 151095818, 168977833}))
  stage_2_butterfly_14 (
    .x_in(stage_1_per_out[28]),
    .y_in(stage_1_per_out[29]),
    .x_out(stage_2_per_in[28]),
    .y_out(stage_2_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({160807241, 177340471, 199876762, 125267062, 260909397, 229100654, 1562592, 55567611,
              43575145, 252241817, 237438985, 42585458, 129101436, 60072008, 1613379, 130696933,
              99187435, 250508912, 77981460, 178386996, 181295312, 64884498, 56094099, 13458851,
              20857483, 27056737, 114486793, 196771169, 61345534, 66242139, 151095818, 168977833}))
  stage_2_butterfly_15 (
    .x_in(stage_1_per_out[30]),
    .y_in(stage_1_per_out[31]),
    .x_out(stage_2_per_in[30]),
    .y_out(stage_2_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({21080194, 126063290, 145034471, 256272276, 44547301, 219083512, 166955734, 237102043,
              218231468, 175719113, 61997323, 156366160, 49504466, 36946189, 11500489, 95861179,
              169480001, 202071175, 34481514, 222683851, 136992892, 225650462, 205961920, 62844488,
              187864761, 266671862, 95282463, 59284831, 5292226, 95560742, 136878682, 138879618}))
  stage_2_butterfly_16 (
    .x_in(stage_1_per_out[32]),
    .y_in(stage_1_per_out[33]),
    .x_out(stage_2_per_in[32]),
    .y_out(stage_2_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({21080194, 126063290, 145034471, 256272276, 44547301, 219083512, 166955734, 237102043,
              218231468, 175719113, 61997323, 156366160, 49504466, 36946189, 11500489, 95861179,
              169480001, 202071175, 34481514, 222683851, 136992892, 225650462, 205961920, 62844488,
              187864761, 266671862, 95282463, 59284831, 5292226, 95560742, 136878682, 138879618}))
  stage_2_butterfly_17 (
    .x_in(stage_1_per_out[34]),
    .y_in(stage_1_per_out[35]),
    .x_out(stage_2_per_in[34]),
    .y_out(stage_2_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({21080194, 126063290, 145034471, 256272276, 44547301, 219083512, 166955734, 237102043,
              218231468, 175719113, 61997323, 156366160, 49504466, 36946189, 11500489, 95861179,
              169480001, 202071175, 34481514, 222683851, 136992892, 225650462, 205961920, 62844488,
              187864761, 266671862, 95282463, 59284831, 5292226, 95560742, 136878682, 138879618}))
  stage_2_butterfly_18 (
    .x_in(stage_1_per_out[36]),
    .y_in(stage_1_per_out[37]),
    .x_out(stage_2_per_in[36]),
    .y_out(stage_2_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({21080194, 126063290, 145034471, 256272276, 44547301, 219083512, 166955734, 237102043,
              218231468, 175719113, 61997323, 156366160, 49504466, 36946189, 11500489, 95861179,
              169480001, 202071175, 34481514, 222683851, 136992892, 225650462, 205961920, 62844488,
              187864761, 266671862, 95282463, 59284831, 5292226, 95560742, 136878682, 138879618}))
  stage_2_butterfly_19 (
    .x_in(stage_1_per_out[38]),
    .y_in(stage_1_per_out[39]),
    .x_out(stage_2_per_in[38]),
    .y_out(stage_2_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({220490426, 97439895, 93740850, 146037274, 58483920, 206649748, 219898221, 10720790,
              251138298, 210914061, 200749611, 143779572, 73698550, 262077011, 242025902, 234350511,
              78649100, 216395023, 263530653, 126520315, 79136411, 224586596, 193296437, 191444307,
              207329882, 243024363, 212214167, 144929841, 58644800, 148390399, 209658551, 206725018}))
  stage_2_butterfly_20 (
    .x_in(stage_1_per_out[40]),
    .y_in(stage_1_per_out[41]),
    .x_out(stage_2_per_in[40]),
    .y_out(stage_2_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({220490426, 97439895, 93740850, 146037274, 58483920, 206649748, 219898221, 10720790,
              251138298, 210914061, 200749611, 143779572, 73698550, 262077011, 242025902, 234350511,
              78649100, 216395023, 263530653, 126520315, 79136411, 224586596, 193296437, 191444307,
              207329882, 243024363, 212214167, 144929841, 58644800, 148390399, 209658551, 206725018}))
  stage_2_butterfly_21 (
    .x_in(stage_1_per_out[42]),
    .y_in(stage_1_per_out[43]),
    .x_out(stage_2_per_in[42]),
    .y_out(stage_2_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({220490426, 97439895, 93740850, 146037274, 58483920, 206649748, 219898221, 10720790,
              251138298, 210914061, 200749611, 143779572, 73698550, 262077011, 242025902, 234350511,
              78649100, 216395023, 263530653, 126520315, 79136411, 224586596, 193296437, 191444307,
              207329882, 243024363, 212214167, 144929841, 58644800, 148390399, 209658551, 206725018}))
  stage_2_butterfly_22 (
    .x_in(stage_1_per_out[44]),
    .y_in(stage_1_per_out[45]),
    .x_out(stage_2_per_in[44]),
    .y_out(stage_2_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({220490426, 97439895, 93740850, 146037274, 58483920, 206649748, 219898221, 10720790,
              251138298, 210914061, 200749611, 143779572, 73698550, 262077011, 242025902, 234350511,
              78649100, 216395023, 263530653, 126520315, 79136411, 224586596, 193296437, 191444307,
              207329882, 243024363, 212214167, 144929841, 58644800, 148390399, 209658551, 206725018}))
  stage_2_butterfly_23 (
    .x_in(stage_1_per_out[46]),
    .y_in(stage_1_per_out[47]),
    .x_out(stage_2_per_in[46]),
    .y_out(stage_2_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({225389748, 164638888, 9810331, 165134943, 74093574, 18298478, 137346680, 10143115,
              154421517, 8950678, 232451599, 225175773, 43078133, 182691070, 247253507, 42156432,
              126188511, 100457939, 24688427, 12196542, 168676526, 234113027, 44301230, 65413984,
              84058929, 113309038, 10003248, 69773246, 68267735, 85252512, 188517169, 140366124}))
  stage_2_butterfly_24 (
    .x_in(stage_1_per_out[48]),
    .y_in(stage_1_per_out[49]),
    .x_out(stage_2_per_in[48]),
    .y_out(stage_2_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({225389748, 164638888, 9810331, 165134943, 74093574, 18298478, 137346680, 10143115,
              154421517, 8950678, 232451599, 225175773, 43078133, 182691070, 247253507, 42156432,
              126188511, 100457939, 24688427, 12196542, 168676526, 234113027, 44301230, 65413984,
              84058929, 113309038, 10003248, 69773246, 68267735, 85252512, 188517169, 140366124}))
  stage_2_butterfly_25 (
    .x_in(stage_1_per_out[50]),
    .y_in(stage_1_per_out[51]),
    .x_out(stage_2_per_in[50]),
    .y_out(stage_2_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({225389748, 164638888, 9810331, 165134943, 74093574, 18298478, 137346680, 10143115,
              154421517, 8950678, 232451599, 225175773, 43078133, 182691070, 247253507, 42156432,
              126188511, 100457939, 24688427, 12196542, 168676526, 234113027, 44301230, 65413984,
              84058929, 113309038, 10003248, 69773246, 68267735, 85252512, 188517169, 140366124}))
  stage_2_butterfly_26 (
    .x_in(stage_1_per_out[52]),
    .y_in(stage_1_per_out[53]),
    .x_out(stage_2_per_in[52]),
    .y_out(stage_2_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({225389748, 164638888, 9810331, 165134943, 74093574, 18298478, 137346680, 10143115,
              154421517, 8950678, 232451599, 225175773, 43078133, 182691070, 247253507, 42156432,
              126188511, 100457939, 24688427, 12196542, 168676526, 234113027, 44301230, 65413984,
              84058929, 113309038, 10003248, 69773246, 68267735, 85252512, 188517169, 140366124}))
  stage_2_butterfly_27 (
    .x_in(stage_1_per_out[54]),
    .y_in(stage_1_per_out[55]),
    .x_out(stage_2_per_in[54]),
    .y_out(stage_2_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({206795535, 10112777, 16471674, 63483304, 64764693, 172935357, 57599709, 66310724,
              40718170, 176665584, 56943278, 171541778, 244216783, 257269778, 232445568, 262358962,
              35754446, 254132077, 219738759, 68736878, 87088032, 5299132, 117221766, 190319963,
              72621624, 85340443, 94612904, 65324949, 57635675, 119568150, 192832423, 73081523}))
  stage_2_butterfly_28 (
    .x_in(stage_1_per_out[56]),
    .y_in(stage_1_per_out[57]),
    .x_out(stage_2_per_in[56]),
    .y_out(stage_2_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({206795535, 10112777, 16471674, 63483304, 64764693, 172935357, 57599709, 66310724,
              40718170, 176665584, 56943278, 171541778, 244216783, 257269778, 232445568, 262358962,
              35754446, 254132077, 219738759, 68736878, 87088032, 5299132, 117221766, 190319963,
              72621624, 85340443, 94612904, 65324949, 57635675, 119568150, 192832423, 73081523}))
  stage_2_butterfly_29 (
    .x_in(stage_1_per_out[58]),
    .y_in(stage_1_per_out[59]),
    .x_out(stage_2_per_in[58]),
    .y_out(stage_2_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({206795535, 10112777, 16471674, 63483304, 64764693, 172935357, 57599709, 66310724,
              40718170, 176665584, 56943278, 171541778, 244216783, 257269778, 232445568, 262358962,
              35754446, 254132077, 219738759, 68736878, 87088032, 5299132, 117221766, 190319963,
              72621624, 85340443, 94612904, 65324949, 57635675, 119568150, 192832423, 73081523}))
  stage_2_butterfly_30 (
    .x_in(stage_1_per_out[60]),
    .y_in(stage_1_per_out[61]),
    .x_out(stage_2_per_in[60]),
    .y_out(stage_2_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({206795535, 10112777, 16471674, 63483304, 64764693, 172935357, 57599709, 66310724,
              40718170, 176665584, 56943278, 171541778, 244216783, 257269778, 232445568, 262358962,
              35754446, 254132077, 219738759, 68736878, 87088032, 5299132, 117221766, 190319963,
              72621624, 85340443, 94612904, 65324949, 57635675, 119568150, 192832423, 73081523}))
  stage_2_butterfly_31 (
    .x_in(stage_1_per_out[62]),
    .y_in(stage_1_per_out[63]),
    .x_out(stage_2_per_in[62]),
    .y_out(stage_2_per_in[63]),
    .clk(clk),
    .rst(rst)
  );




  // TODO(Yang): stage 2 -> stage 3 permutation
  // FIXME: ignore butterfly units for now.
  stage_2_permutation #(
    .DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    .INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_2_3_per (
    .inData_0(stage_2_per_in[0]),
    .inData_1(stage_2_per_in[1]),
    .inData_2(stage_2_per_in[2]),
    .inData_3(stage_2_per_in[3]),
    .inData_4(stage_2_per_in[4]),
    .inData_5(stage_2_per_in[5]),
    .inData_6(stage_2_per_in[6]),
    .inData_7(stage_2_per_in[7]),
    .inData_8(stage_2_per_in[8]),
    .inData_9(stage_2_per_in[9]),
    .inData_10(stage_2_per_in[10]),
    .inData_11(stage_2_per_in[11]),
    .inData_12(stage_2_per_in[12]),
    .inData_13(stage_2_per_in[13]),
    .inData_14(stage_2_per_in[14]),
    .inData_15(stage_2_per_in[15]),
    .inData_16(stage_2_per_in[16]),
    .inData_17(stage_2_per_in[17]),
    .inData_18(stage_2_per_in[18]),
    .inData_19(stage_2_per_in[19]),
    .inData_20(stage_2_per_in[20]),
    .inData_21(stage_2_per_in[21]),
    .inData_22(stage_2_per_in[22]),
    .inData_23(stage_2_per_in[23]),
    .inData_24(stage_2_per_in[24]),
    .inData_25(stage_2_per_in[25]),
    .inData_26(stage_2_per_in[26]),
    .inData_27(stage_2_per_in[27]),
    .inData_28(stage_2_per_in[28]),
    .inData_29(stage_2_per_in[29]),
    .inData_30(stage_2_per_in[30]),
    .inData_31(stage_2_per_in[31]),
    .inData_32(stage_2_per_in[32]),
    .inData_33(stage_2_per_in[33]),
    .inData_34(stage_2_per_in[34]),
    .inData_35(stage_2_per_in[35]),
    .inData_36(stage_2_per_in[36]),
    .inData_37(stage_2_per_in[37]),
    .inData_38(stage_2_per_in[38]),
    .inData_39(stage_2_per_in[39]),
    .inData_40(stage_2_per_in[40]),
    .inData_41(stage_2_per_in[41]),
    .inData_42(stage_2_per_in[42]),
    .inData_43(stage_2_per_in[43]),
    .inData_44(stage_2_per_in[44]),
    .inData_45(stage_2_per_in[45]),
    .inData_46(stage_2_per_in[46]),
    .inData_47(stage_2_per_in[47]),
    .inData_48(stage_2_per_in[48]),
    .inData_49(stage_2_per_in[49]),
    .inData_50(stage_2_per_in[50]),
    .inData_51(stage_2_per_in[51]),
    .inData_52(stage_2_per_in[52]),
    .inData_53(stage_2_per_in[53]),
    .inData_54(stage_2_per_in[54]),
    .inData_55(stage_2_per_in[55]),
    .inData_56(stage_2_per_in[56]),
    .inData_57(stage_2_per_in[57]),
    .inData_58(stage_2_per_in[58]),
    .inData_59(stage_2_per_in[59]),
    .inData_60(stage_2_per_in[60]),
    .inData_61(stage_2_per_in[61]),
    .inData_62(stage_2_per_in[62]),
    .inData_63(stage_2_per_in[63]),
    .outData_0(stage_2_per_out[0]),
    .outData_1(stage_2_per_out[1]),
    .outData_2(stage_2_per_out[2]),
    .outData_3(stage_2_per_out[3]),
    .outData_4(stage_2_per_out[4]),
    .outData_5(stage_2_per_out[5]),
    .outData_6(stage_2_per_out[6]),
    .outData_7(stage_2_per_out[7]),
    .outData_8(stage_2_per_out[8]),
    .outData_9(stage_2_per_out[9]),
    .outData_10(stage_2_per_out[10]),
    .outData_11(stage_2_per_out[11]),
    .outData_12(stage_2_per_out[12]),
    .outData_13(stage_2_per_out[13]),
    .outData_14(stage_2_per_out[14]),
    .outData_15(stage_2_per_out[15]),
    .outData_16(stage_2_per_out[16]),
    .outData_17(stage_2_per_out[17]),
    .outData_18(stage_2_per_out[18]),
    .outData_19(stage_2_per_out[19]),
    .outData_20(stage_2_per_out[20]),
    .outData_21(stage_2_per_out[21]),
    .outData_22(stage_2_per_out[22]),
    .outData_23(stage_2_per_out[23]),
    .outData_24(stage_2_per_out[24]),
    .outData_25(stage_2_per_out[25]),
    .outData_26(stage_2_per_out[26]),
    .outData_27(stage_2_per_out[27]),
    .outData_28(stage_2_per_out[28]),
    .outData_29(stage_2_per_out[29]),
    .outData_30(stage_2_per_out[30]),
    .outData_31(stage_2_per_out[31]),
    .outData_32(stage_2_per_out[32]),
    .outData_33(stage_2_per_out[33]),
    .outData_34(stage_2_per_out[34]),
    .outData_35(stage_2_per_out[35]),
    .outData_36(stage_2_per_out[36]),
    .outData_37(stage_2_per_out[37]),
    .outData_38(stage_2_per_out[38]),
    .outData_39(stage_2_per_out[39]),
    .outData_40(stage_2_per_out[40]),
    .outData_41(stage_2_per_out[41]),
    .outData_42(stage_2_per_out[42]),
    .outData_43(stage_2_per_out[43]),
    .outData_44(stage_2_per_out[44]),
    .outData_45(stage_2_per_out[45]),
    .outData_46(stage_2_per_out[46]),
    .outData_47(stage_2_per_out[47]),
    .outData_48(stage_2_per_out[48]),
    .outData_49(stage_2_per_out[49]),
    .outData_50(stage_2_per_out[50]),
    .outData_51(stage_2_per_out[51]),
    .outData_52(stage_2_per_out[52]),
    .outData_53(stage_2_per_out[53]),
    .outData_54(stage_2_per_out[54]),
    .outData_55(stage_2_per_out[55]),
    .outData_56(stage_2_per_out[56]),
    .outData_57(stage_2_per_out[57]),
    .outData_58(stage_2_per_out[58]),
    .outData_59(stage_2_per_out[59]),
    .outData_60(stage_2_per_out[60]),
    .outData_61(stage_2_per_out[61]),
    .outData_62(stage_2_per_out[62]),
    .outData_63(stage_2_per_out[63]),
    .in_start(in_start[2]),
    .out_start(out_start[2]),
    .clk(clk),
    .rst(rst)
  );

  // TODO(Tian): stage 3 32 butterfly units
  butterfly #(
    .start(START_CYCLE[3]),
    .factors({163812837, 41086336, 77337691, 246744565, 44942358, 63703579, 202221416, 212648666,
              242800442, 210298252, 99962405, 13519489, 98878775, 96648403, 184226747, 22541719,
              186413553, 7055647, 188210893, 71064168, 101839787, 119707826, 170604387, 257798138,
              78777967, 59208162, 91898237, 139182289, 183348420, 9757140, 250166212, 108965460}))
  stage_3_butterfly_0 (
    .x_in(stage_2_per_out[0]),
    .y_in(stage_2_per_out[1]),
    .x_out(stage_3_per_in[0]),
    .y_out(stage_3_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({163812837, 41086336, 77337691, 246744565, 44942358, 63703579, 202221416, 212648666,
              242800442, 210298252, 99962405, 13519489, 98878775, 96648403, 184226747, 22541719,
              186413553, 7055647, 188210893, 71064168, 101839787, 119707826, 170604387, 257798138,
              78777967, 59208162, 91898237, 139182289, 183348420, 9757140, 250166212, 108965460}))
  stage_3_butterfly_1 (
    .x_in(stage_2_per_out[2]),
    .y_in(stage_2_per_out[3]),
    .x_out(stage_3_per_in[2]),
    .y_out(stage_3_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({163812837, 41086336, 77337691, 246744565, 44942358, 63703579, 202221416, 212648666,
              242800442, 210298252, 99962405, 13519489, 98878775, 96648403, 184226747, 22541719,
              186413553, 7055647, 188210893, 71064168, 101839787, 119707826, 170604387, 257798138,
              78777967, 59208162, 91898237, 139182289, 183348420, 9757140, 250166212, 108965460}))
  stage_3_butterfly_2 (
    .x_in(stage_2_per_out[4]),
    .y_in(stage_2_per_out[5]),
    .x_out(stage_3_per_in[4]),
    .y_out(stage_3_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({163812837, 41086336, 77337691, 246744565, 44942358, 63703579, 202221416, 212648666,
              242800442, 210298252, 99962405, 13519489, 98878775, 96648403, 184226747, 22541719,
              186413553, 7055647, 188210893, 71064168, 101839787, 119707826, 170604387, 257798138,
              78777967, 59208162, 91898237, 139182289, 183348420, 9757140, 250166212, 108965460}))
  stage_3_butterfly_3 (
    .x_in(stage_2_per_out[6]),
    .y_in(stage_2_per_out[7]),
    .x_out(stage_3_per_in[6]),
    .y_out(stage_3_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({163812837, 41086336, 77337691, 246744565, 44942358, 63703579, 202221416, 212648666,
              242800442, 210298252, 99962405, 13519489, 98878775, 96648403, 184226747, 22541719,
              186413553, 7055647, 188210893, 71064168, 101839787, 119707826, 170604387, 257798138,
              78777967, 59208162, 91898237, 139182289, 183348420, 9757140, 250166212, 108965460}))
  stage_3_butterfly_4 (
    .x_in(stage_2_per_out[8]),
    .y_in(stage_2_per_out[9]),
    .x_out(stage_3_per_in[8]),
    .y_out(stage_3_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({163812837, 41086336, 77337691, 246744565, 44942358, 63703579, 202221416, 212648666,
              242800442, 210298252, 99962405, 13519489, 98878775, 96648403, 184226747, 22541719,
              186413553, 7055647, 188210893, 71064168, 101839787, 119707826, 170604387, 257798138,
              78777967, 59208162, 91898237, 139182289, 183348420, 9757140, 250166212, 108965460}))
  stage_3_butterfly_5 (
    .x_in(stage_2_per_out[10]),
    .y_in(stage_2_per_out[11]),
    .x_out(stage_3_per_in[10]),
    .y_out(stage_3_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({163812837, 41086336, 77337691, 246744565, 44942358, 63703579, 202221416, 212648666,
              242800442, 210298252, 99962405, 13519489, 98878775, 96648403, 184226747, 22541719,
              186413553, 7055647, 188210893, 71064168, 101839787, 119707826, 170604387, 257798138,
              78777967, 59208162, 91898237, 139182289, 183348420, 9757140, 250166212, 108965460}))
  stage_3_butterfly_6 (
    .x_in(stage_2_per_out[12]),
    .y_in(stage_2_per_out[13]),
    .x_out(stage_3_per_in[12]),
    .y_out(stage_3_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({163812837, 41086336, 77337691, 246744565, 44942358, 63703579, 202221416, 212648666,
              242800442, 210298252, 99962405, 13519489, 98878775, 96648403, 184226747, 22541719,
              186413553, 7055647, 188210893, 71064168, 101839787, 119707826, 170604387, 257798138,
              78777967, 59208162, 91898237, 139182289, 183348420, 9757140, 250166212, 108965460}))
  stage_3_butterfly_7 (
    .x_in(stage_2_per_out[14]),
    .y_in(stage_2_per_out[15]),
    .x_out(stage_3_per_in[14]),
    .y_out(stage_3_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({155168409, 133503098, 34119889, 164195239, 234890903, 241682233, 204152715, 254509489,
              146361539, 197074908, 132703565, 47994339, 258923154, 195631434, 196436059, 13250338,
              176917280, 244883276, 261793746, 101483624, 12328961, 39141691, 13919506, 170227406,
              22463657, 236144340, 83853696, 10130658, 106640438, 59283803, 100484142, 75673633}))
  stage_3_butterfly_8 (
    .x_in(stage_2_per_out[16]),
    .y_in(stage_2_per_out[17]),
    .x_out(stage_3_per_in[16]),
    .y_out(stage_3_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({155168409, 133503098, 34119889, 164195239, 234890903, 241682233, 204152715, 254509489,
              146361539, 197074908, 132703565, 47994339, 258923154, 195631434, 196436059, 13250338,
              176917280, 244883276, 261793746, 101483624, 12328961, 39141691, 13919506, 170227406,
              22463657, 236144340, 83853696, 10130658, 106640438, 59283803, 100484142, 75673633}))
  stage_3_butterfly_9 (
    .x_in(stage_2_per_out[18]),
    .y_in(stage_2_per_out[19]),
    .x_out(stage_3_per_in[18]),
    .y_out(stage_3_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({155168409, 133503098, 34119889, 164195239, 234890903, 241682233, 204152715, 254509489,
              146361539, 197074908, 132703565, 47994339, 258923154, 195631434, 196436059, 13250338,
              176917280, 244883276, 261793746, 101483624, 12328961, 39141691, 13919506, 170227406,
              22463657, 236144340, 83853696, 10130658, 106640438, 59283803, 100484142, 75673633}))
  stage_3_butterfly_10 (
    .x_in(stage_2_per_out[20]),
    .y_in(stage_2_per_out[21]),
    .x_out(stage_3_per_in[20]),
    .y_out(stage_3_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({155168409, 133503098, 34119889, 164195239, 234890903, 241682233, 204152715, 254509489,
              146361539, 197074908, 132703565, 47994339, 258923154, 195631434, 196436059, 13250338,
              176917280, 244883276, 261793746, 101483624, 12328961, 39141691, 13919506, 170227406,
              22463657, 236144340, 83853696, 10130658, 106640438, 59283803, 100484142, 75673633}))
  stage_3_butterfly_11 (
    .x_in(stage_2_per_out[22]),
    .y_in(stage_2_per_out[23]),
    .x_out(stage_3_per_in[22]),
    .y_out(stage_3_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({155168409, 133503098, 34119889, 164195239, 234890903, 241682233, 204152715, 254509489,
              146361539, 197074908, 132703565, 47994339, 258923154, 195631434, 196436059, 13250338,
              176917280, 244883276, 261793746, 101483624, 12328961, 39141691, 13919506, 170227406,
              22463657, 236144340, 83853696, 10130658, 106640438, 59283803, 100484142, 75673633}))
  stage_3_butterfly_12 (
    .x_in(stage_2_per_out[24]),
    .y_in(stage_2_per_out[25]),
    .x_out(stage_3_per_in[24]),
    .y_out(stage_3_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({155168409, 133503098, 34119889, 164195239, 234890903, 241682233, 204152715, 254509489,
              146361539, 197074908, 132703565, 47994339, 258923154, 195631434, 196436059, 13250338,
              176917280, 244883276, 261793746, 101483624, 12328961, 39141691, 13919506, 170227406,
              22463657, 236144340, 83853696, 10130658, 106640438, 59283803, 100484142, 75673633}))
  stage_3_butterfly_13 (
    .x_in(stage_2_per_out[26]),
    .y_in(stage_2_per_out[27]),
    .x_out(stage_3_per_in[26]),
    .y_out(stage_3_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({155168409, 133503098, 34119889, 164195239, 234890903, 241682233, 204152715, 254509489,
              146361539, 197074908, 132703565, 47994339, 258923154, 195631434, 196436059, 13250338,
              176917280, 244883276, 261793746, 101483624, 12328961, 39141691, 13919506, 170227406,
              22463657, 236144340, 83853696, 10130658, 106640438, 59283803, 100484142, 75673633}))
  stage_3_butterfly_14 (
    .x_in(stage_2_per_out[28]),
    .y_in(stage_2_per_out[29]),
    .x_out(stage_3_per_in[28]),
    .y_out(stage_3_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({155168409, 133503098, 34119889, 164195239, 234890903, 241682233, 204152715, 254509489,
              146361539, 197074908, 132703565, 47994339, 258923154, 195631434, 196436059, 13250338,
              176917280, 244883276, 261793746, 101483624, 12328961, 39141691, 13919506, 170227406,
              22463657, 236144340, 83853696, 10130658, 106640438, 59283803, 100484142, 75673633}))
  stage_3_butterfly_15 (
    .x_in(stage_2_per_out[30]),
    .y_in(stage_2_per_out[31]),
    .x_out(stage_3_per_in[30]),
    .y_out(stage_3_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({149528048, 163585105, 201357873, 161827885, 108810259, 40553702, 229216409, 252952333,
              211668928, 147433882, 248876054, 15927889, 28824907, 217644581, 230702770, 69161747,
              189762285, 133081916, 249640399, 257268473, 240677074, 216143425, 123185272, 227894900,
              63350037, 37936257, 241125460, 81777479, 34339674, 173702965, 150873005, 130557622}))
  stage_3_butterfly_16 (
    .x_in(stage_2_per_out[32]),
    .y_in(stage_2_per_out[33]),
    .x_out(stage_3_per_in[32]),
    .y_out(stage_3_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({149528048, 163585105, 201357873, 161827885, 108810259, 40553702, 229216409, 252952333,
              211668928, 147433882, 248876054, 15927889, 28824907, 217644581, 230702770, 69161747,
              189762285, 133081916, 249640399, 257268473, 240677074, 216143425, 123185272, 227894900,
              63350037, 37936257, 241125460, 81777479, 34339674, 173702965, 150873005, 130557622}))
  stage_3_butterfly_17 (
    .x_in(stage_2_per_out[34]),
    .y_in(stage_2_per_out[35]),
    .x_out(stage_3_per_in[34]),
    .y_out(stage_3_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({149528048, 163585105, 201357873, 161827885, 108810259, 40553702, 229216409, 252952333,
              211668928, 147433882, 248876054, 15927889, 28824907, 217644581, 230702770, 69161747,
              189762285, 133081916, 249640399, 257268473, 240677074, 216143425, 123185272, 227894900,
              63350037, 37936257, 241125460, 81777479, 34339674, 173702965, 150873005, 130557622}))
  stage_3_butterfly_18 (
    .x_in(stage_2_per_out[36]),
    .y_in(stage_2_per_out[37]),
    .x_out(stage_3_per_in[36]),
    .y_out(stage_3_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({149528048, 163585105, 201357873, 161827885, 108810259, 40553702, 229216409, 252952333,
              211668928, 147433882, 248876054, 15927889, 28824907, 217644581, 230702770, 69161747,
              189762285, 133081916, 249640399, 257268473, 240677074, 216143425, 123185272, 227894900,
              63350037, 37936257, 241125460, 81777479, 34339674, 173702965, 150873005, 130557622}))
  stage_3_butterfly_19 (
    .x_in(stage_2_per_out[38]),
    .y_in(stage_2_per_out[39]),
    .x_out(stage_3_per_in[38]),
    .y_out(stage_3_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({149528048, 163585105, 201357873, 161827885, 108810259, 40553702, 229216409, 252952333,
              211668928, 147433882, 248876054, 15927889, 28824907, 217644581, 230702770, 69161747,
              189762285, 133081916, 249640399, 257268473, 240677074, 216143425, 123185272, 227894900,
              63350037, 37936257, 241125460, 81777479, 34339674, 173702965, 150873005, 130557622}))
  stage_3_butterfly_20 (
    .x_in(stage_2_per_out[40]),
    .y_in(stage_2_per_out[41]),
    .x_out(stage_3_per_in[40]),
    .y_out(stage_3_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({149528048, 163585105, 201357873, 161827885, 108810259, 40553702, 229216409, 252952333,
              211668928, 147433882, 248876054, 15927889, 28824907, 217644581, 230702770, 69161747,
              189762285, 133081916, 249640399, 257268473, 240677074, 216143425, 123185272, 227894900,
              63350037, 37936257, 241125460, 81777479, 34339674, 173702965, 150873005, 130557622}))
  stage_3_butterfly_21 (
    .x_in(stage_2_per_out[42]),
    .y_in(stage_2_per_out[43]),
    .x_out(stage_3_per_in[42]),
    .y_out(stage_3_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({149528048, 163585105, 201357873, 161827885, 108810259, 40553702, 229216409, 252952333,
              211668928, 147433882, 248876054, 15927889, 28824907, 217644581, 230702770, 69161747,
              189762285, 133081916, 249640399, 257268473, 240677074, 216143425, 123185272, 227894900,
              63350037, 37936257, 241125460, 81777479, 34339674, 173702965, 150873005, 130557622}))
  stage_3_butterfly_22 (
    .x_in(stage_2_per_out[44]),
    .y_in(stage_2_per_out[45]),
    .x_out(stage_3_per_in[44]),
    .y_out(stage_3_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({149528048, 163585105, 201357873, 161827885, 108810259, 40553702, 229216409, 252952333,
              211668928, 147433882, 248876054, 15927889, 28824907, 217644581, 230702770, 69161747,
              189762285, 133081916, 249640399, 257268473, 240677074, 216143425, 123185272, 227894900,
              63350037, 37936257, 241125460, 81777479, 34339674, 173702965, 150873005, 130557622}))
  stage_3_butterfly_23 (
    .x_in(stage_2_per_out[46]),
    .y_in(stage_2_per_out[47]),
    .x_out(stage_3_per_in[46]),
    .y_out(stage_3_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({172227818, 3883583, 41630462, 2795054, 214551729, 149851545, 160286792, 220618744,
              144414946, 42733001, 258649698, 162031725, 139555205, 18399308, 143969713, 87844233,
              246656426, 238498066, 151968102, 68136911, 265950570, 86730411, 85922744, 253827407,
              214085592, 37011073, 25065602, 78488715, 41155851, 90597117, 193371292, 231318087}))
  stage_3_butterfly_24 (
    .x_in(stage_2_per_out[48]),
    .y_in(stage_2_per_out[49]),
    .x_out(stage_3_per_in[48]),
    .y_out(stage_3_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({172227818, 3883583, 41630462, 2795054, 214551729, 149851545, 160286792, 220618744,
              144414946, 42733001, 258649698, 162031725, 139555205, 18399308, 143969713, 87844233,
              246656426, 238498066, 151968102, 68136911, 265950570, 86730411, 85922744, 253827407,
              214085592, 37011073, 25065602, 78488715, 41155851, 90597117, 193371292, 231318087}))
  stage_3_butterfly_25 (
    .x_in(stage_2_per_out[50]),
    .y_in(stage_2_per_out[51]),
    .x_out(stage_3_per_in[50]),
    .y_out(stage_3_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({172227818, 3883583, 41630462, 2795054, 214551729, 149851545, 160286792, 220618744,
              144414946, 42733001, 258649698, 162031725, 139555205, 18399308, 143969713, 87844233,
              246656426, 238498066, 151968102, 68136911, 265950570, 86730411, 85922744, 253827407,
              214085592, 37011073, 25065602, 78488715, 41155851, 90597117, 193371292, 231318087}))
  stage_3_butterfly_26 (
    .x_in(stage_2_per_out[52]),
    .y_in(stage_2_per_out[53]),
    .x_out(stage_3_per_in[52]),
    .y_out(stage_3_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({172227818, 3883583, 41630462, 2795054, 214551729, 149851545, 160286792, 220618744,
              144414946, 42733001, 258649698, 162031725, 139555205, 18399308, 143969713, 87844233,
              246656426, 238498066, 151968102, 68136911, 265950570, 86730411, 85922744, 253827407,
              214085592, 37011073, 25065602, 78488715, 41155851, 90597117, 193371292, 231318087}))
  stage_3_butterfly_27 (
    .x_in(stage_2_per_out[54]),
    .y_in(stage_2_per_out[55]),
    .x_out(stage_3_per_in[54]),
    .y_out(stage_3_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({172227818, 3883583, 41630462, 2795054, 214551729, 149851545, 160286792, 220618744,
              144414946, 42733001, 258649698, 162031725, 139555205, 18399308, 143969713, 87844233,
              246656426, 238498066, 151968102, 68136911, 265950570, 86730411, 85922744, 253827407,
              214085592, 37011073, 25065602, 78488715, 41155851, 90597117, 193371292, 231318087}))
  stage_3_butterfly_28 (
    .x_in(stage_2_per_out[56]),
    .y_in(stage_2_per_out[57]),
    .x_out(stage_3_per_in[56]),
    .y_out(stage_3_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({172227818, 3883583, 41630462, 2795054, 214551729, 149851545, 160286792, 220618744,
              144414946, 42733001, 258649698, 162031725, 139555205, 18399308, 143969713, 87844233,
              246656426, 238498066, 151968102, 68136911, 265950570, 86730411, 85922744, 253827407,
              214085592, 37011073, 25065602, 78488715, 41155851, 90597117, 193371292, 231318087}))
  stage_3_butterfly_29 (
    .x_in(stage_2_per_out[58]),
    .y_in(stage_2_per_out[59]),
    .x_out(stage_3_per_in[58]),
    .y_out(stage_3_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({172227818, 3883583, 41630462, 2795054, 214551729, 149851545, 160286792, 220618744,
              144414946, 42733001, 258649698, 162031725, 139555205, 18399308, 143969713, 87844233,
              246656426, 238498066, 151968102, 68136911, 265950570, 86730411, 85922744, 253827407,
              214085592, 37011073, 25065602, 78488715, 41155851, 90597117, 193371292, 231318087}))
  stage_3_butterfly_30 (
    .x_in(stage_2_per_out[60]),
    .y_in(stage_2_per_out[61]),
    .x_out(stage_3_per_in[60]),
    .y_out(stage_3_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({172227818, 3883583, 41630462, 2795054, 214551729, 149851545, 160286792, 220618744,
              144414946, 42733001, 258649698, 162031725, 139555205, 18399308, 143969713, 87844233,
              246656426, 238498066, 151968102, 68136911, 265950570, 86730411, 85922744, 253827407,
              214085592, 37011073, 25065602, 78488715, 41155851, 90597117, 193371292, 231318087}))
  stage_3_butterfly_31 (
    .x_in(stage_2_per_out[62]),
    .y_in(stage_2_per_out[63]),
    .x_out(stage_3_per_in[62]),
    .y_out(stage_3_per_in[63]),
    .clk(clk),
    .rst(rst)
  );



  // TODO(Yang): stage 3 -> stage 4 permutation
  // FIXME: ignore butterfly units for now.
  stage_3_permutation #(
    .DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    .INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_3_4_per (
    .inData_0(stage_3_per_in[0]),
    .inData_1(stage_3_per_in[1]),
    .inData_2(stage_3_per_in[2]),
    .inData_3(stage_3_per_in[3]),
    .inData_4(stage_3_per_in[4]),
    .inData_5(stage_3_per_in[5]),
    .inData_6(stage_3_per_in[6]),
    .inData_7(stage_3_per_in[7]),
    .inData_8(stage_3_per_in[8]),
    .inData_9(stage_3_per_in[9]),
    .inData_10(stage_3_per_in[10]),
    .inData_11(stage_3_per_in[11]),
    .inData_12(stage_3_per_in[12]),
    .inData_13(stage_3_per_in[13]),
    .inData_14(stage_3_per_in[14]),
    .inData_15(stage_3_per_in[15]),
    .inData_16(stage_3_per_in[16]),
    .inData_17(stage_3_per_in[17]),
    .inData_18(stage_3_per_in[18]),
    .inData_19(stage_3_per_in[19]),
    .inData_20(stage_3_per_in[20]),
    .inData_21(stage_3_per_in[21]),
    .inData_22(stage_3_per_in[22]),
    .inData_23(stage_3_per_in[23]),
    .inData_24(stage_3_per_in[24]),
    .inData_25(stage_3_per_in[25]),
    .inData_26(stage_3_per_in[26]),
    .inData_27(stage_3_per_in[27]),
    .inData_28(stage_3_per_in[28]),
    .inData_29(stage_3_per_in[29]),
    .inData_30(stage_3_per_in[30]),
    .inData_31(stage_3_per_in[31]),
    .inData_32(stage_3_per_in[32]),
    .inData_33(stage_3_per_in[33]),
    .inData_34(stage_3_per_in[34]),
    .inData_35(stage_3_per_in[35]),
    .inData_36(stage_3_per_in[36]),
    .inData_37(stage_3_per_in[37]),
    .inData_38(stage_3_per_in[38]),
    .inData_39(stage_3_per_in[39]),
    .inData_40(stage_3_per_in[40]),
    .inData_41(stage_3_per_in[41]),
    .inData_42(stage_3_per_in[42]),
    .inData_43(stage_3_per_in[43]),
    .inData_44(stage_3_per_in[44]),
    .inData_45(stage_3_per_in[45]),
    .inData_46(stage_3_per_in[46]),
    .inData_47(stage_3_per_in[47]),
    .inData_48(stage_3_per_in[48]),
    .inData_49(stage_3_per_in[49]),
    .inData_50(stage_3_per_in[50]),
    .inData_51(stage_3_per_in[51]),
    .inData_52(stage_3_per_in[52]),
    .inData_53(stage_3_per_in[53]),
    .inData_54(stage_3_per_in[54]),
    .inData_55(stage_3_per_in[55]),
    .inData_56(stage_3_per_in[56]),
    .inData_57(stage_3_per_in[57]),
    .inData_58(stage_3_per_in[58]),
    .inData_59(stage_3_per_in[59]),
    .inData_60(stage_3_per_in[60]),
    .inData_61(stage_3_per_in[61]),
    .inData_62(stage_3_per_in[62]),
    .inData_63(stage_3_per_in[63]),
    .outData_0(stage_3_per_out[0]),
    .outData_1(stage_3_per_out[1]),
    .outData_2(stage_3_per_out[2]),
    .outData_3(stage_3_per_out[3]),
    .outData_4(stage_3_per_out[4]),
    .outData_5(stage_3_per_out[5]),
    .outData_6(stage_3_per_out[6]),
    .outData_7(stage_3_per_out[7]),
    .outData_8(stage_3_per_out[8]),
    .outData_9(stage_3_per_out[9]),
    .outData_10(stage_3_per_out[10]),
    .outData_11(stage_3_per_out[11]),
    .outData_12(stage_3_per_out[12]),
    .outData_13(stage_3_per_out[13]),
    .outData_14(stage_3_per_out[14]),
    .outData_15(stage_3_per_out[15]),
    .outData_16(stage_3_per_out[16]),
    .outData_17(stage_3_per_out[17]),
    .outData_18(stage_3_per_out[18]),
    .outData_19(stage_3_per_out[19]),
    .outData_20(stage_3_per_out[20]),
    .outData_21(stage_3_per_out[21]),
    .outData_22(stage_3_per_out[22]),
    .outData_23(stage_3_per_out[23]),
    .outData_24(stage_3_per_out[24]),
    .outData_25(stage_3_per_out[25]),
    .outData_26(stage_3_per_out[26]),
    .outData_27(stage_3_per_out[27]),
    .outData_28(stage_3_per_out[28]),
    .outData_29(stage_3_per_out[29]),
    .outData_30(stage_3_per_out[30]),
    .outData_31(stage_3_per_out[31]),
    .outData_32(stage_3_per_out[32]),
    .outData_33(stage_3_per_out[33]),
    .outData_34(stage_3_per_out[34]),
    .outData_35(stage_3_per_out[35]),
    .outData_36(stage_3_per_out[36]),
    .outData_37(stage_3_per_out[37]),
    .outData_38(stage_3_per_out[38]),
    .outData_39(stage_3_per_out[39]),
    .outData_40(stage_3_per_out[40]),
    .outData_41(stage_3_per_out[41]),
    .outData_42(stage_3_per_out[42]),
    .outData_43(stage_3_per_out[43]),
    .outData_44(stage_3_per_out[44]),
    .outData_45(stage_3_per_out[45]),
    .outData_46(stage_3_per_out[46]),
    .outData_47(stage_3_per_out[47]),
    .outData_48(stage_3_per_out[48]),
    .outData_49(stage_3_per_out[49]),
    .outData_50(stage_3_per_out[50]),
    .outData_51(stage_3_per_out[51]),
    .outData_52(stage_3_per_out[52]),
    .outData_53(stage_3_per_out[53]),
    .outData_54(stage_3_per_out[54]),
    .outData_55(stage_3_per_out[55]),
    .outData_56(stage_3_per_out[56]),
    .outData_57(stage_3_per_out[57]),
    .outData_58(stage_3_per_out[58]),
    .outData_59(stage_3_per_out[59]),
    .outData_60(stage_3_per_out[60]),
    .outData_61(stage_3_per_out[61]),
    .outData_62(stage_3_per_out[62]),
    .outData_63(stage_3_per_out[63]),
    .in_start(in_start[3]),
    .out_start(out_start[3]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 4 32 butterfly units
  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 215696667, 153962078, 233560477, 181852808, 146694818, 218546733, 227611463,
              17079898, 25574347, 263678998, 27685019, 179817683, 6323336, 200054106, 170752771,
              141548072, 70982951, 124918999, 39593842, 102065274, 109254766, 237620966, 210568560,
              76642651, 201062854, 152865265, 62045777, 168270865, 235204060, 162373432, 112472991}))
  stage_4_butterfly_0 (
    .x_in(stage_3_per_out[0]),
    .y_in(stage_3_per_out[1]),
    .x_out(stage_4_per_in[0]),
    .y_out(stage_4_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 215696667, 153962078, 233560477, 181852808, 146694818, 218546733, 227611463,
              17079898, 25574347, 263678998, 27685019, 179817683, 6323336, 200054106, 170752771,
              141548072, 70982951, 124918999, 39593842, 102065274, 109254766, 237620966, 210568560,
              76642651, 201062854, 152865265, 62045777, 168270865, 235204060, 162373432, 112472991}))
  stage_4_butterfly_1 (
    .x_in(stage_3_per_out[2]),
    .y_in(stage_3_per_out[3]),
    .x_out(stage_4_per_in[2]),
    .y_out(stage_4_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 215696667, 153962078, 233560477, 181852808, 146694818, 218546733, 227611463,
              17079898, 25574347, 263678998, 27685019, 179817683, 6323336, 200054106, 170752771,
              141548072, 70982951, 124918999, 39593842, 102065274, 109254766, 237620966, 210568560,
              76642651, 201062854, 152865265, 62045777, 168270865, 235204060, 162373432, 112472991}))
  stage_4_butterfly_2 (
    .x_in(stage_3_per_out[4]),
    .y_in(stage_3_per_out[5]),
    .x_out(stage_4_per_in[4]),
    .y_out(stage_4_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 215696667, 153962078, 233560477, 181852808, 146694818, 218546733, 227611463,
              17079898, 25574347, 263678998, 27685019, 179817683, 6323336, 200054106, 170752771,
              141548072, 70982951, 124918999, 39593842, 102065274, 109254766, 237620966, 210568560,
              76642651, 201062854, 152865265, 62045777, 168270865, 235204060, 162373432, 112472991}))
  stage_4_butterfly_3 (
    .x_in(stage_3_per_out[6]),
    .y_in(stage_3_per_out[7]),
    .x_out(stage_4_per_in[6]),
    .y_out(stage_4_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 215696667, 153962078, 233560477, 181852808, 146694818, 218546733, 227611463,
              17079898, 25574347, 263678998, 27685019, 179817683, 6323336, 200054106, 170752771,
              141548072, 70982951, 124918999, 39593842, 102065274, 109254766, 237620966, 210568560,
              76642651, 201062854, 152865265, 62045777, 168270865, 235204060, 162373432, 112472991}))
  stage_4_butterfly_4 (
    .x_in(stage_3_per_out[8]),
    .y_in(stage_3_per_out[9]),
    .x_out(stage_4_per_in[8]),
    .y_out(stage_4_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 215696667, 153962078, 233560477, 181852808, 146694818, 218546733, 227611463,
              17079898, 25574347, 263678998, 27685019, 179817683, 6323336, 200054106, 170752771,
              141548072, 70982951, 124918999, 39593842, 102065274, 109254766, 237620966, 210568560,
              76642651, 201062854, 152865265, 62045777, 168270865, 235204060, 162373432, 112472991}))
  stage_4_butterfly_5 (
    .x_in(stage_3_per_out[10]),
    .y_in(stage_3_per_out[11]),
    .x_out(stage_4_per_in[10]),
    .y_out(stage_4_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 215696667, 153962078, 233560477, 181852808, 146694818, 218546733, 227611463,
              17079898, 25574347, 263678998, 27685019, 179817683, 6323336, 200054106, 170752771,
              141548072, 70982951, 124918999, 39593842, 102065274, 109254766, 237620966, 210568560,
              76642651, 201062854, 152865265, 62045777, 168270865, 235204060, 162373432, 112472991}))
  stage_4_butterfly_6 (
    .x_in(stage_3_per_out[12]),
    .y_in(stage_3_per_out[13]),
    .x_out(stage_4_per_in[12]),
    .y_out(stage_4_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 215696667, 153962078, 233560477, 181852808, 146694818, 218546733, 227611463,
              17079898, 25574347, 263678998, 27685019, 179817683, 6323336, 200054106, 170752771,
              141548072, 70982951, 124918999, 39593842, 102065274, 109254766, 237620966, 210568560,
              76642651, 201062854, 152865265, 62045777, 168270865, 235204060, 162373432, 112472991}))
  stage_4_butterfly_7 (
    .x_in(stage_3_per_out[14]),
    .y_in(stage_3_per_out[15]),
    .x_out(stage_4_per_in[14]),
    .y_out(stage_4_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 215696667, 153962078, 233560477, 181852808, 146694818, 218546733, 227611463,
              17079898, 25574347, 263678998, 27685019, 179817683, 6323336, 200054106, 170752771,
              141548072, 70982951, 124918999, 39593842, 102065274, 109254766, 237620966, 210568560,
              76642651, 201062854, 152865265, 62045777, 168270865, 235204060, 162373432, 112472991}))
  stage_4_butterfly_8 (
    .x_in(stage_3_per_out[16]),
    .y_in(stage_3_per_out[17]),
    .x_out(stage_4_per_in[16]),
    .y_out(stage_4_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 215696667, 153962078, 233560477, 181852808, 146694818, 218546733, 227611463,
              17079898, 25574347, 263678998, 27685019, 179817683, 6323336, 200054106, 170752771,
              141548072, 70982951, 124918999, 39593842, 102065274, 109254766, 237620966, 210568560,
              76642651, 201062854, 152865265, 62045777, 168270865, 235204060, 162373432, 112472991}))
  stage_4_butterfly_9 (
    .x_in(stage_3_per_out[18]),
    .y_in(stage_3_per_out[19]),
    .x_out(stage_4_per_in[18]),
    .y_out(stage_4_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 215696667, 153962078, 233560477, 181852808, 146694818, 218546733, 227611463,
              17079898, 25574347, 263678998, 27685019, 179817683, 6323336, 200054106, 170752771,
              141548072, 70982951, 124918999, 39593842, 102065274, 109254766, 237620966, 210568560,
              76642651, 201062854, 152865265, 62045777, 168270865, 235204060, 162373432, 112472991}))
  stage_4_butterfly_10 (
    .x_in(stage_3_per_out[20]),
    .y_in(stage_3_per_out[21]),
    .x_out(stage_4_per_in[20]),
    .y_out(stage_4_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 215696667, 153962078, 233560477, 181852808, 146694818, 218546733, 227611463,
              17079898, 25574347, 263678998, 27685019, 179817683, 6323336, 200054106, 170752771,
              141548072, 70982951, 124918999, 39593842, 102065274, 109254766, 237620966, 210568560,
              76642651, 201062854, 152865265, 62045777, 168270865, 235204060, 162373432, 112472991}))
  stage_4_butterfly_11 (
    .x_in(stage_3_per_out[22]),
    .y_in(stage_3_per_out[23]),
    .x_out(stage_4_per_in[22]),
    .y_out(stage_4_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 215696667, 153962078, 233560477, 181852808, 146694818, 218546733, 227611463,
              17079898, 25574347, 263678998, 27685019, 179817683, 6323336, 200054106, 170752771,
              141548072, 70982951, 124918999, 39593842, 102065274, 109254766, 237620966, 210568560,
              76642651, 201062854, 152865265, 62045777, 168270865, 235204060, 162373432, 112472991}))
  stage_4_butterfly_12 (
    .x_in(stage_3_per_out[24]),
    .y_in(stage_3_per_out[25]),
    .x_out(stage_4_per_in[24]),
    .y_out(stage_4_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 215696667, 153962078, 233560477, 181852808, 146694818, 218546733, 227611463,
              17079898, 25574347, 263678998, 27685019, 179817683, 6323336, 200054106, 170752771,
              141548072, 70982951, 124918999, 39593842, 102065274, 109254766, 237620966, 210568560,
              76642651, 201062854, 152865265, 62045777, 168270865, 235204060, 162373432, 112472991}))
  stage_4_butterfly_13 (
    .x_in(stage_3_per_out[26]),
    .y_in(stage_3_per_out[27]),
    .x_out(stage_4_per_in[26]),
    .y_out(stage_4_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 215696667, 153962078, 233560477, 181852808, 146694818, 218546733, 227611463,
              17079898, 25574347, 263678998, 27685019, 179817683, 6323336, 200054106, 170752771,
              141548072, 70982951, 124918999, 39593842, 102065274, 109254766, 237620966, 210568560,
              76642651, 201062854, 152865265, 62045777, 168270865, 235204060, 162373432, 112472991}))
  stage_4_butterfly_14 (
    .x_in(stage_3_per_out[28]),
    .y_in(stage_3_per_out[29]),
    .x_out(stage_4_per_in[28]),
    .y_out(stage_4_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 215696667, 153962078, 233560477, 181852808, 146694818, 218546733, 227611463,
              17079898, 25574347, 263678998, 27685019, 179817683, 6323336, 200054106, 170752771,
              141548072, 70982951, 124918999, 39593842, 102065274, 109254766, 237620966, 210568560,
              76642651, 201062854, 152865265, 62045777, 168270865, 235204060, 162373432, 112472991}))
  stage_4_butterfly_15 (
    .x_in(stage_3_per_out[30]),
    .y_in(stage_3_per_out[31]),
    .x_out(stage_4_per_in[30]),
    .y_out(stage_4_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({197787791, 172642311, 11695616, 189907315, 147699054, 202366126, 78852289, 71460019,
              193045667, 66112528, 115957373, 47317233, 109553202, 165226744, 191662816, 140204941,
              169276669, 119224607, 82771912, 239095400, 157085730, 208403048, 111341228, 177255039,
              41084242, 130295133, 175609590, 118939950, 71471012, 131798756, 74680748, 145384235}))
  stage_4_butterfly_16 (
    .x_in(stage_3_per_out[32]),
    .y_in(stage_3_per_out[33]),
    .x_out(stage_4_per_in[32]),
    .y_out(stage_4_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({197787791, 172642311, 11695616, 189907315, 147699054, 202366126, 78852289, 71460019,
              193045667, 66112528, 115957373, 47317233, 109553202, 165226744, 191662816, 140204941,
              169276669, 119224607, 82771912, 239095400, 157085730, 208403048, 111341228, 177255039,
              41084242, 130295133, 175609590, 118939950, 71471012, 131798756, 74680748, 145384235}))
  stage_4_butterfly_17 (
    .x_in(stage_3_per_out[34]),
    .y_in(stage_3_per_out[35]),
    .x_out(stage_4_per_in[34]),
    .y_out(stage_4_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({197787791, 172642311, 11695616, 189907315, 147699054, 202366126, 78852289, 71460019,
              193045667, 66112528, 115957373, 47317233, 109553202, 165226744, 191662816, 140204941,
              169276669, 119224607, 82771912, 239095400, 157085730, 208403048, 111341228, 177255039,
              41084242, 130295133, 175609590, 118939950, 71471012, 131798756, 74680748, 145384235}))
  stage_4_butterfly_18 (
    .x_in(stage_3_per_out[36]),
    .y_in(stage_3_per_out[37]),
    .x_out(stage_4_per_in[36]),
    .y_out(stage_4_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({197787791, 172642311, 11695616, 189907315, 147699054, 202366126, 78852289, 71460019,
              193045667, 66112528, 115957373, 47317233, 109553202, 165226744, 191662816, 140204941,
              169276669, 119224607, 82771912, 239095400, 157085730, 208403048, 111341228, 177255039,
              41084242, 130295133, 175609590, 118939950, 71471012, 131798756, 74680748, 145384235}))
  stage_4_butterfly_19 (
    .x_in(stage_3_per_out[38]),
    .y_in(stage_3_per_out[39]),
    .x_out(stage_4_per_in[38]),
    .y_out(stage_4_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({197787791, 172642311, 11695616, 189907315, 147699054, 202366126, 78852289, 71460019,
              193045667, 66112528, 115957373, 47317233, 109553202, 165226744, 191662816, 140204941,
              169276669, 119224607, 82771912, 239095400, 157085730, 208403048, 111341228, 177255039,
              41084242, 130295133, 175609590, 118939950, 71471012, 131798756, 74680748, 145384235}))
  stage_4_butterfly_20 (
    .x_in(stage_3_per_out[40]),
    .y_in(stage_3_per_out[41]),
    .x_out(stage_4_per_in[40]),
    .y_out(stage_4_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({197787791, 172642311, 11695616, 189907315, 147699054, 202366126, 78852289, 71460019,
              193045667, 66112528, 115957373, 47317233, 109553202, 165226744, 191662816, 140204941,
              169276669, 119224607, 82771912, 239095400, 157085730, 208403048, 111341228, 177255039,
              41084242, 130295133, 175609590, 118939950, 71471012, 131798756, 74680748, 145384235}))
  stage_4_butterfly_21 (
    .x_in(stage_3_per_out[42]),
    .y_in(stage_3_per_out[43]),
    .x_out(stage_4_per_in[42]),
    .y_out(stage_4_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({197787791, 172642311, 11695616, 189907315, 147699054, 202366126, 78852289, 71460019,
              193045667, 66112528, 115957373, 47317233, 109553202, 165226744, 191662816, 140204941,
              169276669, 119224607, 82771912, 239095400, 157085730, 208403048, 111341228, 177255039,
              41084242, 130295133, 175609590, 118939950, 71471012, 131798756, 74680748, 145384235}))
  stage_4_butterfly_22 (
    .x_in(stage_3_per_out[44]),
    .y_in(stage_3_per_out[45]),
    .x_out(stage_4_per_in[44]),
    .y_out(stage_4_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({197787791, 172642311, 11695616, 189907315, 147699054, 202366126, 78852289, 71460019,
              193045667, 66112528, 115957373, 47317233, 109553202, 165226744, 191662816, 140204941,
              169276669, 119224607, 82771912, 239095400, 157085730, 208403048, 111341228, 177255039,
              41084242, 130295133, 175609590, 118939950, 71471012, 131798756, 74680748, 145384235}))
  stage_4_butterfly_23 (
    .x_in(stage_3_per_out[46]),
    .y_in(stage_3_per_out[47]),
    .x_out(stage_4_per_in[46]),
    .y_out(stage_4_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({197787791, 172642311, 11695616, 189907315, 147699054, 202366126, 78852289, 71460019,
              193045667, 66112528, 115957373, 47317233, 109553202, 165226744, 191662816, 140204941,
              169276669, 119224607, 82771912, 239095400, 157085730, 208403048, 111341228, 177255039,
              41084242, 130295133, 175609590, 118939950, 71471012, 131798756, 74680748, 145384235}))
  stage_4_butterfly_24 (
    .x_in(stage_3_per_out[48]),
    .y_in(stage_3_per_out[49]),
    .x_out(stage_4_per_in[48]),
    .y_out(stage_4_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({197787791, 172642311, 11695616, 189907315, 147699054, 202366126, 78852289, 71460019,
              193045667, 66112528, 115957373, 47317233, 109553202, 165226744, 191662816, 140204941,
              169276669, 119224607, 82771912, 239095400, 157085730, 208403048, 111341228, 177255039,
              41084242, 130295133, 175609590, 118939950, 71471012, 131798756, 74680748, 145384235}))
  stage_4_butterfly_25 (
    .x_in(stage_3_per_out[50]),
    .y_in(stage_3_per_out[51]),
    .x_out(stage_4_per_in[50]),
    .y_out(stage_4_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({197787791, 172642311, 11695616, 189907315, 147699054, 202366126, 78852289, 71460019,
              193045667, 66112528, 115957373, 47317233, 109553202, 165226744, 191662816, 140204941,
              169276669, 119224607, 82771912, 239095400, 157085730, 208403048, 111341228, 177255039,
              41084242, 130295133, 175609590, 118939950, 71471012, 131798756, 74680748, 145384235}))
  stage_4_butterfly_26 (
    .x_in(stage_3_per_out[52]),
    .y_in(stage_3_per_out[53]),
    .x_out(stage_4_per_in[52]),
    .y_out(stage_4_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({197787791, 172642311, 11695616, 189907315, 147699054, 202366126, 78852289, 71460019,
              193045667, 66112528, 115957373, 47317233, 109553202, 165226744, 191662816, 140204941,
              169276669, 119224607, 82771912, 239095400, 157085730, 208403048, 111341228, 177255039,
              41084242, 130295133, 175609590, 118939950, 71471012, 131798756, 74680748, 145384235}))
  stage_4_butterfly_27 (
    .x_in(stage_3_per_out[54]),
    .y_in(stage_3_per_out[55]),
    .x_out(stage_4_per_in[54]),
    .y_out(stage_4_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({197787791, 172642311, 11695616, 189907315, 147699054, 202366126, 78852289, 71460019,
              193045667, 66112528, 115957373, 47317233, 109553202, 165226744, 191662816, 140204941,
              169276669, 119224607, 82771912, 239095400, 157085730, 208403048, 111341228, 177255039,
              41084242, 130295133, 175609590, 118939950, 71471012, 131798756, 74680748, 145384235}))
  stage_4_butterfly_28 (
    .x_in(stage_3_per_out[56]),
    .y_in(stage_3_per_out[57]),
    .x_out(stage_4_per_in[56]),
    .y_out(stage_4_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({197787791, 172642311, 11695616, 189907315, 147699054, 202366126, 78852289, 71460019,
              193045667, 66112528, 115957373, 47317233, 109553202, 165226744, 191662816, 140204941,
              169276669, 119224607, 82771912, 239095400, 157085730, 208403048, 111341228, 177255039,
              41084242, 130295133, 175609590, 118939950, 71471012, 131798756, 74680748, 145384235}))
  stage_4_butterfly_29 (
    .x_in(stage_3_per_out[58]),
    .y_in(stage_3_per_out[59]),
    .x_out(stage_4_per_in[58]),
    .y_out(stage_4_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({197787791, 172642311, 11695616, 189907315, 147699054, 202366126, 78852289, 71460019,
              193045667, 66112528, 115957373, 47317233, 109553202, 165226744, 191662816, 140204941,
              169276669, 119224607, 82771912, 239095400, 157085730, 208403048, 111341228, 177255039,
              41084242, 130295133, 175609590, 118939950, 71471012, 131798756, 74680748, 145384235}))
  stage_4_butterfly_30 (
    .x_in(stage_3_per_out[60]),
    .y_in(stage_3_per_out[61]),
    .x_out(stage_4_per_in[60]),
    .y_out(stage_4_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({197787791, 172642311, 11695616, 189907315, 147699054, 202366126, 78852289, 71460019,
              193045667, 66112528, 115957373, 47317233, 109553202, 165226744, 191662816, 140204941,
              169276669, 119224607, 82771912, 239095400, 157085730, 208403048, 111341228, 177255039,
              41084242, 130295133, 175609590, 118939950, 71471012, 131798756, 74680748, 145384235}))
  stage_4_butterfly_31 (
    .x_in(stage_3_per_out[62]),
    .y_in(stage_3_per_out[63]),
    .x_out(stage_4_per_in[62]),
    .y_out(stage_4_per_in[63]),
    .clk(clk),
    .rst(rst)
  );



  // TODO(Yang): stage 4 -> stage 5 permutation
  // FIXME: ignore butterfly units for now.
  stage_4_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_4_5_per (
    .inData_0(stage_4_per_in[0]),
    .inData_1(stage_4_per_in[1]),
    .inData_2(stage_4_per_in[2]),
    .inData_3(stage_4_per_in[3]),
    .inData_4(stage_4_per_in[4]),
    .inData_5(stage_4_per_in[5]),
    .inData_6(stage_4_per_in[6]),
    .inData_7(stage_4_per_in[7]),
    .inData_8(stage_4_per_in[8]),
    .inData_9(stage_4_per_in[9]),
    .inData_10(stage_4_per_in[10]),
    .inData_11(stage_4_per_in[11]),
    .inData_12(stage_4_per_in[12]),
    .inData_13(stage_4_per_in[13]),
    .inData_14(stage_4_per_in[14]),
    .inData_15(stage_4_per_in[15]),
    .inData_16(stage_4_per_in[16]),
    .inData_17(stage_4_per_in[17]),
    .inData_18(stage_4_per_in[18]),
    .inData_19(stage_4_per_in[19]),
    .inData_20(stage_4_per_in[20]),
    .inData_21(stage_4_per_in[21]),
    .inData_22(stage_4_per_in[22]),
    .inData_23(stage_4_per_in[23]),
    .inData_24(stage_4_per_in[24]),
    .inData_25(stage_4_per_in[25]),
    .inData_26(stage_4_per_in[26]),
    .inData_27(stage_4_per_in[27]),
    .inData_28(stage_4_per_in[28]),
    .inData_29(stage_4_per_in[29]),
    .inData_30(stage_4_per_in[30]),
    .inData_31(stage_4_per_in[31]),
    .inData_32(stage_4_per_in[32]),
    .inData_33(stage_4_per_in[33]),
    .inData_34(stage_4_per_in[34]),
    .inData_35(stage_4_per_in[35]),
    .inData_36(stage_4_per_in[36]),
    .inData_37(stage_4_per_in[37]),
    .inData_38(stage_4_per_in[38]),
    .inData_39(stage_4_per_in[39]),
    .inData_40(stage_4_per_in[40]),
    .inData_41(stage_4_per_in[41]),
    .inData_42(stage_4_per_in[42]),
    .inData_43(stage_4_per_in[43]),
    .inData_44(stage_4_per_in[44]),
    .inData_45(stage_4_per_in[45]),
    .inData_46(stage_4_per_in[46]),
    .inData_47(stage_4_per_in[47]),
    .inData_48(stage_4_per_in[48]),
    .inData_49(stage_4_per_in[49]),
    .inData_50(stage_4_per_in[50]),
    .inData_51(stage_4_per_in[51]),
    .inData_52(stage_4_per_in[52]),
    .inData_53(stage_4_per_in[53]),
    .inData_54(stage_4_per_in[54]),
    .inData_55(stage_4_per_in[55]),
    .inData_56(stage_4_per_in[56]),
    .inData_57(stage_4_per_in[57]),
    .inData_58(stage_4_per_in[58]),
    .inData_59(stage_4_per_in[59]),
    .inData_60(stage_4_per_in[60]),
    .inData_61(stage_4_per_in[61]),
    .inData_62(stage_4_per_in[62]),
    .inData_63(stage_4_per_in[63]),
    .outData_0(stage_4_per_out[0]),
    .outData_1(stage_4_per_out[1]),
    .outData_2(stage_4_per_out[2]),
    .outData_3(stage_4_per_out[3]),
    .outData_4(stage_4_per_out[4]),
    .outData_5(stage_4_per_out[5]),
    .outData_6(stage_4_per_out[6]),
    .outData_7(stage_4_per_out[7]),
    .outData_8(stage_4_per_out[8]),
    .outData_9(stage_4_per_out[9]),
    .outData_10(stage_4_per_out[10]),
    .outData_11(stage_4_per_out[11]),
    .outData_12(stage_4_per_out[12]),
    .outData_13(stage_4_per_out[13]),
    .outData_14(stage_4_per_out[14]),
    .outData_15(stage_4_per_out[15]),
    .outData_16(stage_4_per_out[16]),
    .outData_17(stage_4_per_out[17]),
    .outData_18(stage_4_per_out[18]),
    .outData_19(stage_4_per_out[19]),
    .outData_20(stage_4_per_out[20]),
    .outData_21(stage_4_per_out[21]),
    .outData_22(stage_4_per_out[22]),
    .outData_23(stage_4_per_out[23]),
    .outData_24(stage_4_per_out[24]),
    .outData_25(stage_4_per_out[25]),
    .outData_26(stage_4_per_out[26]),
    .outData_27(stage_4_per_out[27]),
    .outData_28(stage_4_per_out[28]),
    .outData_29(stage_4_per_out[29]),
    .outData_30(stage_4_per_out[30]),
    .outData_31(stage_4_per_out[31]),
    .outData_32(stage_4_per_out[32]),
    .outData_33(stage_4_per_out[33]),
    .outData_34(stage_4_per_out[34]),
    .outData_35(stage_4_per_out[35]),
    .outData_36(stage_4_per_out[36]),
    .outData_37(stage_4_per_out[37]),
    .outData_38(stage_4_per_out[38]),
    .outData_39(stage_4_per_out[39]),
    .outData_40(stage_4_per_out[40]),
    .outData_41(stage_4_per_out[41]),
    .outData_42(stage_4_per_out[42]),
    .outData_43(stage_4_per_out[43]),
    .outData_44(stage_4_per_out[44]),
    .outData_45(stage_4_per_out[45]),
    .outData_46(stage_4_per_out[46]),
    .outData_47(stage_4_per_out[47]),
    .outData_48(stage_4_per_out[48]),
    .outData_49(stage_4_per_out[49]),
    .outData_50(stage_4_per_out[50]),
    .outData_51(stage_4_per_out[51]),
    .outData_52(stage_4_per_out[52]),
    .outData_53(stage_4_per_out[53]),
    .outData_54(stage_4_per_out[54]),
    .outData_55(stage_4_per_out[55]),
    .outData_56(stage_4_per_out[56]),
    .outData_57(stage_4_per_out[57]),
    .outData_58(stage_4_per_out[58]),
    .outData_59(stage_4_per_out[59]),
    .outData_60(stage_4_per_out[60]),
    .outData_61(stage_4_per_out[61]),
    .outData_62(stage_4_per_out[62]),
    .outData_63(stage_4_per_out[63]),
    .in_start(in_start[4]),
    .out_start(out_start[4]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 5 32 butterfly units
  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_0 (
    .x_in(stage_4_per_out[0]),
    .y_in(stage_4_per_out[1]),
    .x_out(stage_5_per_in[0]),
    .y_out(stage_5_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_1 (
    .x_in(stage_4_per_out[2]),
    .y_in(stage_4_per_out[3]),
    .x_out(stage_5_per_in[2]),
    .y_out(stage_5_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_2 (
    .x_in(stage_4_per_out[4]),
    .y_in(stage_4_per_out[5]),
    .x_out(stage_5_per_in[4]),
    .y_out(stage_5_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_3 (
    .x_in(stage_4_per_out[6]),
    .y_in(stage_4_per_out[7]),
    .x_out(stage_5_per_in[6]),
    .y_out(stage_5_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_4 (
    .x_in(stage_4_per_out[8]),
    .y_in(stage_4_per_out[9]),
    .x_out(stage_5_per_in[8]),
    .y_out(stage_5_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_5 (
    .x_in(stage_4_per_out[10]),
    .y_in(stage_4_per_out[11]),
    .x_out(stage_5_per_in[10]),
    .y_out(stage_5_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_6 (
    .x_in(stage_4_per_out[12]),
    .y_in(stage_4_per_out[13]),
    .x_out(stage_5_per_in[12]),
    .y_out(stage_5_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_7 (
    .x_in(stage_4_per_out[14]),
    .y_in(stage_4_per_out[15]),
    .x_out(stage_5_per_in[14]),
    .y_out(stage_5_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_8 (
    .x_in(stage_4_per_out[16]),
    .y_in(stage_4_per_out[17]),
    .x_out(stage_5_per_in[16]),
    .y_out(stage_5_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_9 (
    .x_in(stage_4_per_out[18]),
    .y_in(stage_4_per_out[19]),
    .x_out(stage_5_per_in[18]),
    .y_out(stage_5_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_10 (
    .x_in(stage_4_per_out[20]),
    .y_in(stage_4_per_out[21]),
    .x_out(stage_5_per_in[20]),
    .y_out(stage_5_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_11 (
    .x_in(stage_4_per_out[22]),
    .y_in(stage_4_per_out[23]),
    .x_out(stage_5_per_in[22]),
    .y_out(stage_5_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_12 (
    .x_in(stage_4_per_out[24]),
    .y_in(stage_4_per_out[25]),
    .x_out(stage_5_per_in[24]),
    .y_out(stage_5_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_13 (
    .x_in(stage_4_per_out[26]),
    .y_in(stage_4_per_out[27]),
    .x_out(stage_5_per_in[26]),
    .y_out(stage_5_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_14 (
    .x_in(stage_4_per_out[28]),
    .y_in(stage_4_per_out[29]),
    .x_out(stage_5_per_in[28]),
    .y_out(stage_5_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_15 (
    .x_in(stage_4_per_out[30]),
    .y_in(stage_4_per_out[31]),
    .x_out(stage_5_per_in[30]),
    .y_out(stage_5_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_16 (
    .x_in(stage_4_per_out[32]),
    .y_in(stage_4_per_out[33]),
    .x_out(stage_5_per_in[32]),
    .y_out(stage_5_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_17 (
    .x_in(stage_4_per_out[34]),
    .y_in(stage_4_per_out[35]),
    .x_out(stage_5_per_in[34]),
    .y_out(stage_5_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_18 (
    .x_in(stage_4_per_out[36]),
    .y_in(stage_4_per_out[37]),
    .x_out(stage_5_per_in[36]),
    .y_out(stage_5_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_19 (
    .x_in(stage_4_per_out[38]),
    .y_in(stage_4_per_out[39]),
    .x_out(stage_5_per_in[38]),
    .y_out(stage_5_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_20 (
    .x_in(stage_4_per_out[40]),
    .y_in(stage_4_per_out[41]),
    .x_out(stage_5_per_in[40]),
    .y_out(stage_5_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_21 (
    .x_in(stage_4_per_out[42]),
    .y_in(stage_4_per_out[43]),
    .x_out(stage_5_per_in[42]),
    .y_out(stage_5_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_22 (
    .x_in(stage_4_per_out[44]),
    .y_in(stage_4_per_out[45]),
    .x_out(stage_5_per_in[44]),
    .y_out(stage_5_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_23 (
    .x_in(stage_4_per_out[46]),
    .y_in(stage_4_per_out[47]),
    .x_out(stage_5_per_in[46]),
    .y_out(stage_5_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_24 (
    .x_in(stage_4_per_out[48]),
    .y_in(stage_4_per_out[49]),
    .x_out(stage_5_per_in[48]),
    .y_out(stage_5_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_25 (
    .x_in(stage_4_per_out[50]),
    .y_in(stage_4_per_out[51]),
    .x_out(stage_5_per_in[50]),
    .y_out(stage_5_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_26 (
    .x_in(stage_4_per_out[52]),
    .y_in(stage_4_per_out[53]),
    .x_out(stage_5_per_in[52]),
    .y_out(stage_5_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_27 (
    .x_in(stage_4_per_out[54]),
    .y_in(stage_4_per_out[55]),
    .x_out(stage_5_per_in[54]),
    .y_out(stage_5_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_28 (
    .x_in(stage_4_per_out[56]),
    .y_in(stage_4_per_out[57]),
    .x_out(stage_5_per_in[56]),
    .y_out(stage_5_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_29 (
    .x_in(stage_4_per_out[58]),
    .y_in(stage_4_per_out[59]),
    .x_out(stage_5_per_in[58]),
    .y_out(stage_5_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_30 (
    .x_in(stage_4_per_out[60]),
    .y_in(stage_4_per_out[61]),
    .x_out(stage_5_per_in[60]),
    .y_out(stage_5_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 108349160, 178374402, 220656190, 174234737, 36955649, 216372172, 221840088,
              249274747, 206308099, 35289455, 76573097, 11699091, 143639106, 234642902, 39264098,
              57538295, 84893967, 265190919, 165596304, 102579498, 119480423, 139368110, 72061017,
              92744225, 5258704, 83571649, 220492738, 18533839, 99790517, 196317032, 73825164}))
  stage_5_butterfly_31 (
    .x_in(stage_4_per_out[62]),
    .y_in(stage_4_per_out[63]),
    .x_out(stage_5_per_in[62]),
    .y_out(stage_5_per_in[63]),
    .clk(clk),
    .rst(rst)
  );



  // TODO(Yang): stage 5 -> stage 6 permutation
  // FIXME: ignore butterfly units for now.
  stage_5_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_5_6_per (
    .inData_0(stage_5_per_in[0]),
    .inData_1(stage_5_per_in[1]),
    .inData_2(stage_5_per_in[2]),
    .inData_3(stage_5_per_in[3]),
    .inData_4(stage_5_per_in[4]),
    .inData_5(stage_5_per_in[5]),
    .inData_6(stage_5_per_in[6]),
    .inData_7(stage_5_per_in[7]),
    .inData_8(stage_5_per_in[8]),
    .inData_9(stage_5_per_in[9]),
    .inData_10(stage_5_per_in[10]),
    .inData_11(stage_5_per_in[11]),
    .inData_12(stage_5_per_in[12]),
    .inData_13(stage_5_per_in[13]),
    .inData_14(stage_5_per_in[14]),
    .inData_15(stage_5_per_in[15]),
    .inData_16(stage_5_per_in[16]),
    .inData_17(stage_5_per_in[17]),
    .inData_18(stage_5_per_in[18]),
    .inData_19(stage_5_per_in[19]),
    .inData_20(stage_5_per_in[20]),
    .inData_21(stage_5_per_in[21]),
    .inData_22(stage_5_per_in[22]),
    .inData_23(stage_5_per_in[23]),
    .inData_24(stage_5_per_in[24]),
    .inData_25(stage_5_per_in[25]),
    .inData_26(stage_5_per_in[26]),
    .inData_27(stage_5_per_in[27]),
    .inData_28(stage_5_per_in[28]),
    .inData_29(stage_5_per_in[29]),
    .inData_30(stage_5_per_in[30]),
    .inData_31(stage_5_per_in[31]),
    .inData_32(stage_5_per_in[32]),
    .inData_33(stage_5_per_in[33]),
    .inData_34(stage_5_per_in[34]),
    .inData_35(stage_5_per_in[35]),
    .inData_36(stage_5_per_in[36]),
    .inData_37(stage_5_per_in[37]),
    .inData_38(stage_5_per_in[38]),
    .inData_39(stage_5_per_in[39]),
    .inData_40(stage_5_per_in[40]),
    .inData_41(stage_5_per_in[41]),
    .inData_42(stage_5_per_in[42]),
    .inData_43(stage_5_per_in[43]),
    .inData_44(stage_5_per_in[44]),
    .inData_45(stage_5_per_in[45]),
    .inData_46(stage_5_per_in[46]),
    .inData_47(stage_5_per_in[47]),
    .inData_48(stage_5_per_in[48]),
    .inData_49(stage_5_per_in[49]),
    .inData_50(stage_5_per_in[50]),
    .inData_51(stage_5_per_in[51]),
    .inData_52(stage_5_per_in[52]),
    .inData_53(stage_5_per_in[53]),
    .inData_54(stage_5_per_in[54]),
    .inData_55(stage_5_per_in[55]),
    .inData_56(stage_5_per_in[56]),
    .inData_57(stage_5_per_in[57]),
    .inData_58(stage_5_per_in[58]),
    .inData_59(stage_5_per_in[59]),
    .inData_60(stage_5_per_in[60]),
    .inData_61(stage_5_per_in[61]),
    .inData_62(stage_5_per_in[62]),
    .inData_63(stage_5_per_in[63]),
    .outData_0(stage_5_per_out[0]),
    .outData_1(stage_5_per_out[1]),
    .outData_2(stage_5_per_out[2]),
    .outData_3(stage_5_per_out[3]),
    .outData_4(stage_5_per_out[4]),
    .outData_5(stage_5_per_out[5]),
    .outData_6(stage_5_per_out[6]),
    .outData_7(stage_5_per_out[7]),
    .outData_8(stage_5_per_out[8]),
    .outData_9(stage_5_per_out[9]),
    .outData_10(stage_5_per_out[10]),
    .outData_11(stage_5_per_out[11]),
    .outData_12(stage_5_per_out[12]),
    .outData_13(stage_5_per_out[13]),
    .outData_14(stage_5_per_out[14]),
    .outData_15(stage_5_per_out[15]),
    .outData_16(stage_5_per_out[16]),
    .outData_17(stage_5_per_out[17]),
    .outData_18(stage_5_per_out[18]),
    .outData_19(stage_5_per_out[19]),
    .outData_20(stage_5_per_out[20]),
    .outData_21(stage_5_per_out[21]),
    .outData_22(stage_5_per_out[22]),
    .outData_23(stage_5_per_out[23]),
    .outData_24(stage_5_per_out[24]),
    .outData_25(stage_5_per_out[25]),
    .outData_26(stage_5_per_out[26]),
    .outData_27(stage_5_per_out[27]),
    .outData_28(stage_5_per_out[28]),
    .outData_29(stage_5_per_out[29]),
    .outData_30(stage_5_per_out[30]),
    .outData_31(stage_5_per_out[31]),
    .outData_32(stage_5_per_out[32]),
    .outData_33(stage_5_per_out[33]),
    .outData_34(stage_5_per_out[34]),
    .outData_35(stage_5_per_out[35]),
    .outData_36(stage_5_per_out[36]),
    .outData_37(stage_5_per_out[37]),
    .outData_38(stage_5_per_out[38]),
    .outData_39(stage_5_per_out[39]),
    .outData_40(stage_5_per_out[40]),
    .outData_41(stage_5_per_out[41]),
    .outData_42(stage_5_per_out[42]),
    .outData_43(stage_5_per_out[43]),
    .outData_44(stage_5_per_out[44]),
    .outData_45(stage_5_per_out[45]),
    .outData_46(stage_5_per_out[46]),
    .outData_47(stage_5_per_out[47]),
    .outData_48(stage_5_per_out[48]),
    .outData_49(stage_5_per_out[49]),
    .outData_50(stage_5_per_out[50]),
    .outData_51(stage_5_per_out[51]),
    .outData_52(stage_5_per_out[52]),
    .outData_53(stage_5_per_out[53]),
    .outData_54(stage_5_per_out[54]),
    .outData_55(stage_5_per_out[55]),
    .outData_56(stage_5_per_out[56]),
    .outData_57(stage_5_per_out[57]),
    .outData_58(stage_5_per_out[58]),
    .outData_59(stage_5_per_out[59]),
    .outData_60(stage_5_per_out[60]),
    .outData_61(stage_5_per_out[61]),
    .outData_62(stage_5_per_out[62]),
    .outData_63(stage_5_per_out[63]),
    .in_start(in_start[5]),
    .out_start(out_start[5]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 6 32 butterfly units
  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_0 (
    .x_in(stage_5_per_out[0]),
    .y_in(stage_5_per_out[1]),
    .x_out(stage_6_per_in[0]),
    .y_out(stage_6_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_1 (
    .x_in(stage_5_per_out[2]),
    .y_in(stage_5_per_out[3]),
    .x_out(stage_6_per_in[2]),
    .y_out(stage_6_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_2 (
    .x_in(stage_5_per_out[4]),
    .y_in(stage_5_per_out[5]),
    .x_out(stage_6_per_in[4]),
    .y_out(stage_6_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_3 (
    .x_in(stage_5_per_out[6]),
    .y_in(stage_5_per_out[7]),
    .x_out(stage_6_per_in[6]),
    .y_out(stage_6_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_4 (
    .x_in(stage_5_per_out[8]),
    .y_in(stage_5_per_out[9]),
    .x_out(stage_6_per_in[8]),
    .y_out(stage_6_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_5 (
    .x_in(stage_5_per_out[10]),
    .y_in(stage_5_per_out[11]),
    .x_out(stage_6_per_in[10]),
    .y_out(stage_6_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_6 (
    .x_in(stage_5_per_out[12]),
    .y_in(stage_5_per_out[13]),
    .x_out(stage_6_per_in[12]),
    .y_out(stage_6_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_7 (
    .x_in(stage_5_per_out[14]),
    .y_in(stage_5_per_out[15]),
    .x_out(stage_6_per_in[14]),
    .y_out(stage_6_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_8 (
    .x_in(stage_5_per_out[16]),
    .y_in(stage_5_per_out[17]),
    .x_out(stage_6_per_in[16]),
    .y_out(stage_6_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_9 (
    .x_in(stage_5_per_out[18]),
    .y_in(stage_5_per_out[19]),
    .x_out(stage_6_per_in[18]),
    .y_out(stage_6_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_10 (
    .x_in(stage_5_per_out[20]),
    .y_in(stage_5_per_out[21]),
    .x_out(stage_6_per_in[20]),
    .y_out(stage_6_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_11 (
    .x_in(stage_5_per_out[22]),
    .y_in(stage_5_per_out[23]),
    .x_out(stage_6_per_in[22]),
    .y_out(stage_6_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_12 (
    .x_in(stage_5_per_out[24]),
    .y_in(stage_5_per_out[25]),
    .x_out(stage_6_per_in[24]),
    .y_out(stage_6_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_13 (
    .x_in(stage_5_per_out[26]),
    .y_in(stage_5_per_out[27]),
    .x_out(stage_6_per_in[26]),
    .y_out(stage_6_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_14 (
    .x_in(stage_5_per_out[28]),
    .y_in(stage_5_per_out[29]),
    .x_out(stage_6_per_in[28]),
    .y_out(stage_6_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_15 (
    .x_in(stage_5_per_out[30]),
    .y_in(stage_5_per_out[31]),
    .x_out(stage_6_per_in[30]),
    .y_out(stage_6_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_16 (
    .x_in(stage_5_per_out[32]),
    .y_in(stage_5_per_out[33]),
    .x_out(stage_6_per_in[32]),
    .y_out(stage_6_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_17 (
    .x_in(stage_5_per_out[34]),
    .y_in(stage_5_per_out[35]),
    .x_out(stage_6_per_in[34]),
    .y_out(stage_6_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_18 (
    .x_in(stage_5_per_out[36]),
    .y_in(stage_5_per_out[37]),
    .x_out(stage_6_per_in[36]),
    .y_out(stage_6_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_19 (
    .x_in(stage_5_per_out[38]),
    .y_in(stage_5_per_out[39]),
    .x_out(stage_6_per_in[38]),
    .y_out(stage_6_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_20 (
    .x_in(stage_5_per_out[40]),
    .y_in(stage_5_per_out[41]),
    .x_out(stage_6_per_in[40]),
    .y_out(stage_6_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_21 (
    .x_in(stage_5_per_out[42]),
    .y_in(stage_5_per_out[43]),
    .x_out(stage_6_per_in[42]),
    .y_out(stage_6_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_22 (
    .x_in(stage_5_per_out[44]),
    .y_in(stage_5_per_out[45]),
    .x_out(stage_6_per_in[44]),
    .y_out(stage_6_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_23 (
    .x_in(stage_5_per_out[46]),
    .y_in(stage_5_per_out[47]),
    .x_out(stage_6_per_in[46]),
    .y_out(stage_6_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_24 (
    .x_in(stage_5_per_out[48]),
    .y_in(stage_5_per_out[49]),
    .x_out(stage_6_per_in[48]),
    .y_out(stage_6_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_25 (
    .x_in(stage_5_per_out[50]),
    .y_in(stage_5_per_out[51]),
    .x_out(stage_6_per_in[50]),
    .y_out(stage_6_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_26 (
    .x_in(stage_5_per_out[52]),
    .y_in(stage_5_per_out[53]),
    .x_out(stage_6_per_in[52]),
    .y_out(stage_6_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_27 (
    .x_in(stage_5_per_out[54]),
    .y_in(stage_5_per_out[55]),
    .x_out(stage_6_per_in[54]),
    .y_out(stage_6_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_28 (
    .x_in(stage_5_per_out[56]),
    .y_in(stage_5_per_out[57]),
    .x_out(stage_6_per_in[56]),
    .y_out(stage_6_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_29 (
    .x_in(stage_5_per_out[58]),
    .y_in(stage_5_per_out[59]),
    .x_out(stage_6_per_in[58]),
    .y_out(stage_6_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_30 (
    .x_in(stage_5_per_out[60]),
    .y_in(stage_5_per_out[61]),
    .x_out(stage_6_per_in[60]),
    .y_out(stage_6_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 163057267, 163057267, 42982065, 42982065, 135333989, 135333989,
              46265048, 46265048, 242569099, 242569099, 70516281, 70516281, 136955445, 136955445,
              33383981, 33383981, 47600907, 47600907, 142393906, 142393906, 69075086, 69075086,
              210749829, 210749829, 133782759, 133782759, 155624840, 155624840, 7802111, 7802111}))
  stage_6_butterfly_31 (
    .x_in(stage_5_per_out[62]),
    .y_in(stage_5_per_out[63]),
    .x_out(stage_6_per_in[62]),
    .y_out(stage_6_per_in[63]),
    .clk(clk),
    .rst(rst)
  );



  // TODO(Yang): stage 6 -> stage 7 permutation
  // FIXME: ignore butterfly units for now.
  stage_6_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_6_7_per (
    .inData_0(stage_6_per_in[0]),
    .inData_1(stage_6_per_in[1]),
    .inData_2(stage_6_per_in[2]),
    .inData_3(stage_6_per_in[3]),
    .inData_4(stage_6_per_in[4]),
    .inData_5(stage_6_per_in[5]),
    .inData_6(stage_6_per_in[6]),
    .inData_7(stage_6_per_in[7]),
    .inData_8(stage_6_per_in[8]),
    .inData_9(stage_6_per_in[9]),
    .inData_10(stage_6_per_in[10]),
    .inData_11(stage_6_per_in[11]),
    .inData_12(stage_6_per_in[12]),
    .inData_13(stage_6_per_in[13]),
    .inData_14(stage_6_per_in[14]),
    .inData_15(stage_6_per_in[15]),
    .inData_16(stage_6_per_in[16]),
    .inData_17(stage_6_per_in[17]),
    .inData_18(stage_6_per_in[18]),
    .inData_19(stage_6_per_in[19]),
    .inData_20(stage_6_per_in[20]),
    .inData_21(stage_6_per_in[21]),
    .inData_22(stage_6_per_in[22]),
    .inData_23(stage_6_per_in[23]),
    .inData_24(stage_6_per_in[24]),
    .inData_25(stage_6_per_in[25]),
    .inData_26(stage_6_per_in[26]),
    .inData_27(stage_6_per_in[27]),
    .inData_28(stage_6_per_in[28]),
    .inData_29(stage_6_per_in[29]),
    .inData_30(stage_6_per_in[30]),
    .inData_31(stage_6_per_in[31]),
    .inData_32(stage_6_per_in[32]),
    .inData_33(stage_6_per_in[33]),
    .inData_34(stage_6_per_in[34]),
    .inData_35(stage_6_per_in[35]),
    .inData_36(stage_6_per_in[36]),
    .inData_37(stage_6_per_in[37]),
    .inData_38(stage_6_per_in[38]),
    .inData_39(stage_6_per_in[39]),
    .inData_40(stage_6_per_in[40]),
    .inData_41(stage_6_per_in[41]),
    .inData_42(stage_6_per_in[42]),
    .inData_43(stage_6_per_in[43]),
    .inData_44(stage_6_per_in[44]),
    .inData_45(stage_6_per_in[45]),
    .inData_46(stage_6_per_in[46]),
    .inData_47(stage_6_per_in[47]),
    .inData_48(stage_6_per_in[48]),
    .inData_49(stage_6_per_in[49]),
    .inData_50(stage_6_per_in[50]),
    .inData_51(stage_6_per_in[51]),
    .inData_52(stage_6_per_in[52]),
    .inData_53(stage_6_per_in[53]),
    .inData_54(stage_6_per_in[54]),
    .inData_55(stage_6_per_in[55]),
    .inData_56(stage_6_per_in[56]),
    .inData_57(stage_6_per_in[57]),
    .inData_58(stage_6_per_in[58]),
    .inData_59(stage_6_per_in[59]),
    .inData_60(stage_6_per_in[60]),
    .inData_61(stage_6_per_in[61]),
    .inData_62(stage_6_per_in[62]),
    .inData_63(stage_6_per_in[63]),
    .outData_0(stage_6_per_out[0]),
    .outData_1(stage_6_per_out[1]),
    .outData_2(stage_6_per_out[2]),
    .outData_3(stage_6_per_out[3]),
    .outData_4(stage_6_per_out[4]),
    .outData_5(stage_6_per_out[5]),
    .outData_6(stage_6_per_out[6]),
    .outData_7(stage_6_per_out[7]),
    .outData_8(stage_6_per_out[8]),
    .outData_9(stage_6_per_out[9]),
    .outData_10(stage_6_per_out[10]),
    .outData_11(stage_6_per_out[11]),
    .outData_12(stage_6_per_out[12]),
    .outData_13(stage_6_per_out[13]),
    .outData_14(stage_6_per_out[14]),
    .outData_15(stage_6_per_out[15]),
    .outData_16(stage_6_per_out[16]),
    .outData_17(stage_6_per_out[17]),
    .outData_18(stage_6_per_out[18]),
    .outData_19(stage_6_per_out[19]),
    .outData_20(stage_6_per_out[20]),
    .outData_21(stage_6_per_out[21]),
    .outData_22(stage_6_per_out[22]),
    .outData_23(stage_6_per_out[23]),
    .outData_24(stage_6_per_out[24]),
    .outData_25(stage_6_per_out[25]),
    .outData_26(stage_6_per_out[26]),
    .outData_27(stage_6_per_out[27]),
    .outData_28(stage_6_per_out[28]),
    .outData_29(stage_6_per_out[29]),
    .outData_30(stage_6_per_out[30]),
    .outData_31(stage_6_per_out[31]),
    .outData_32(stage_6_per_out[32]),
    .outData_33(stage_6_per_out[33]),
    .outData_34(stage_6_per_out[34]),
    .outData_35(stage_6_per_out[35]),
    .outData_36(stage_6_per_out[36]),
    .outData_37(stage_6_per_out[37]),
    .outData_38(stage_6_per_out[38]),
    .outData_39(stage_6_per_out[39]),
    .outData_40(stage_6_per_out[40]),
    .outData_41(stage_6_per_out[41]),
    .outData_42(stage_6_per_out[42]),
    .outData_43(stage_6_per_out[43]),
    .outData_44(stage_6_per_out[44]),
    .outData_45(stage_6_per_out[45]),
    .outData_46(stage_6_per_out[46]),
    .outData_47(stage_6_per_out[47]),
    .outData_48(stage_6_per_out[48]),
    .outData_49(stage_6_per_out[49]),
    .outData_50(stage_6_per_out[50]),
    .outData_51(stage_6_per_out[51]),
    .outData_52(stage_6_per_out[52]),
    .outData_53(stage_6_per_out[53]),
    .outData_54(stage_6_per_out[54]),
    .outData_55(stage_6_per_out[55]),
    .outData_56(stage_6_per_out[56]),
    .outData_57(stage_6_per_out[57]),
    .outData_58(stage_6_per_out[58]),
    .outData_59(stage_6_per_out[59]),
    .outData_60(stage_6_per_out[60]),
    .outData_61(stage_6_per_out[61]),
    .outData_62(stage_6_per_out[62]),
    .outData_63(stage_6_per_out[63]),
    .in_start(in_start[6]),
    .out_start(out_start[6]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 7 32 butterfly units
  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_0 (
    .x_in(stage_6_per_out[0]),
    .y_in(stage_6_per_out[1]),
    .x_out(stage_7_per_in[0]),
    .y_out(stage_7_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_1 (
    .x_in(stage_6_per_out[2]),
    .y_in(stage_6_per_out[3]),
    .x_out(stage_7_per_in[2]),
    .y_out(stage_7_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_2 (
    .x_in(stage_6_per_out[4]),
    .y_in(stage_6_per_out[5]),
    .x_out(stage_7_per_in[4]),
    .y_out(stage_7_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_3 (
    .x_in(stage_6_per_out[6]),
    .y_in(stage_6_per_out[7]),
    .x_out(stage_7_per_in[6]),
    .y_out(stage_7_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_4 (
    .x_in(stage_6_per_out[8]),
    .y_in(stage_6_per_out[9]),
    .x_out(stage_7_per_in[8]),
    .y_out(stage_7_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_5 (
    .x_in(stage_6_per_out[10]),
    .y_in(stage_6_per_out[11]),
    .x_out(stage_7_per_in[10]),
    .y_out(stage_7_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_6 (
    .x_in(stage_6_per_out[12]),
    .y_in(stage_6_per_out[13]),
    .x_out(stage_7_per_in[12]),
    .y_out(stage_7_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_7 (
    .x_in(stage_6_per_out[14]),
    .y_in(stage_6_per_out[15]),
    .x_out(stage_7_per_in[14]),
    .y_out(stage_7_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_8 (
    .x_in(stage_6_per_out[16]),
    .y_in(stage_6_per_out[17]),
    .x_out(stage_7_per_in[16]),
    .y_out(stage_7_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_9 (
    .x_in(stage_6_per_out[18]),
    .y_in(stage_6_per_out[19]),
    .x_out(stage_7_per_in[18]),
    .y_out(stage_7_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_10 (
    .x_in(stage_6_per_out[20]),
    .y_in(stage_6_per_out[21]),
    .x_out(stage_7_per_in[20]),
    .y_out(stage_7_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_11 (
    .x_in(stage_6_per_out[22]),
    .y_in(stage_6_per_out[23]),
    .x_out(stage_7_per_in[22]),
    .y_out(stage_7_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_12 (
    .x_in(stage_6_per_out[24]),
    .y_in(stage_6_per_out[25]),
    .x_out(stage_7_per_in[24]),
    .y_out(stage_7_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_13 (
    .x_in(stage_6_per_out[26]),
    .y_in(stage_6_per_out[27]),
    .x_out(stage_7_per_in[26]),
    .y_out(stage_7_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_14 (
    .x_in(stage_6_per_out[28]),
    .y_in(stage_6_per_out[29]),
    .x_out(stage_7_per_in[28]),
    .y_out(stage_7_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_15 (
    .x_in(stage_6_per_out[30]),
    .y_in(stage_6_per_out[31]),
    .x_out(stage_7_per_in[30]),
    .y_out(stage_7_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_16 (
    .x_in(stage_6_per_out[32]),
    .y_in(stage_6_per_out[33]),
    .x_out(stage_7_per_in[32]),
    .y_out(stage_7_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_17 (
    .x_in(stage_6_per_out[34]),
    .y_in(stage_6_per_out[35]),
    .x_out(stage_7_per_in[34]),
    .y_out(stage_7_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_18 (
    .x_in(stage_6_per_out[36]),
    .y_in(stage_6_per_out[37]),
    .x_out(stage_7_per_in[36]),
    .y_out(stage_7_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_19 (
    .x_in(stage_6_per_out[38]),
    .y_in(stage_6_per_out[39]),
    .x_out(stage_7_per_in[38]),
    .y_out(stage_7_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_20 (
    .x_in(stage_6_per_out[40]),
    .y_in(stage_6_per_out[41]),
    .x_out(stage_7_per_in[40]),
    .y_out(stage_7_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_21 (
    .x_in(stage_6_per_out[42]),
    .y_in(stage_6_per_out[43]),
    .x_out(stage_7_per_in[42]),
    .y_out(stage_7_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_22 (
    .x_in(stage_6_per_out[44]),
    .y_in(stage_6_per_out[45]),
    .x_out(stage_7_per_in[44]),
    .y_out(stage_7_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_23 (
    .x_in(stage_6_per_out[46]),
    .y_in(stage_6_per_out[47]),
    .x_out(stage_7_per_in[46]),
    .y_out(stage_7_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_24 (
    .x_in(stage_6_per_out[48]),
    .y_in(stage_6_per_out[49]),
    .x_out(stage_7_per_in[48]),
    .y_out(stage_7_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_25 (
    .x_in(stage_6_per_out[50]),
    .y_in(stage_6_per_out[51]),
    .x_out(stage_7_per_in[50]),
    .y_out(stage_7_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_26 (
    .x_in(stage_6_per_out[52]),
    .y_in(stage_6_per_out[53]),
    .x_out(stage_7_per_in[52]),
    .y_out(stage_7_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_27 (
    .x_in(stage_6_per_out[54]),
    .y_in(stage_6_per_out[55]),
    .x_out(stage_7_per_in[54]),
    .y_out(stage_7_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_28 (
    .x_in(stage_6_per_out[56]),
    .y_in(stage_6_per_out[57]),
    .x_out(stage_7_per_in[56]),
    .y_out(stage_7_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_29 (
    .x_in(stage_6_per_out[58]),
    .y_in(stage_6_per_out[59]),
    .x_out(stage_7_per_in[58]),
    .y_out(stage_7_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_30 (
    .x_in(stage_6_per_out[60]),
    .y_in(stage_6_per_out[61]),
    .x_out(stage_7_per_in[60]),
    .y_out(stage_7_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_31 (
    .x_in(stage_6_per_out[62]),
    .y_in(stage_6_per_out[63]),
    .x_out(stage_7_per_in[62]),
    .y_out(stage_7_per_in[63]),
    .clk(clk),
    .rst(rst)
  );



  // TODO(Yang): stage 7 -> stage 8 permutation
  // FIXME: ignore butterfly units for now.
  stage_7_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_7_8_per (
    .inData_0(stage_7_per_in[0]),
    .inData_1(stage_7_per_in[1]),
    .inData_2(stage_7_per_in[2]),
    .inData_3(stage_7_per_in[3]),
    .inData_4(stage_7_per_in[4]),
    .inData_5(stage_7_per_in[5]),
    .inData_6(stage_7_per_in[6]),
    .inData_7(stage_7_per_in[7]),
    .inData_8(stage_7_per_in[8]),
    .inData_9(stage_7_per_in[9]),
    .inData_10(stage_7_per_in[10]),
    .inData_11(stage_7_per_in[11]),
    .inData_12(stage_7_per_in[12]),
    .inData_13(stage_7_per_in[13]),
    .inData_14(stage_7_per_in[14]),
    .inData_15(stage_7_per_in[15]),
    .inData_16(stage_7_per_in[16]),
    .inData_17(stage_7_per_in[17]),
    .inData_18(stage_7_per_in[18]),
    .inData_19(stage_7_per_in[19]),
    .inData_20(stage_7_per_in[20]),
    .inData_21(stage_7_per_in[21]),
    .inData_22(stage_7_per_in[22]),
    .inData_23(stage_7_per_in[23]),
    .inData_24(stage_7_per_in[24]),
    .inData_25(stage_7_per_in[25]),
    .inData_26(stage_7_per_in[26]),
    .inData_27(stage_7_per_in[27]),
    .inData_28(stage_7_per_in[28]),
    .inData_29(stage_7_per_in[29]),
    .inData_30(stage_7_per_in[30]),
    .inData_31(stage_7_per_in[31]),
    .inData_32(stage_7_per_in[32]),
    .inData_33(stage_7_per_in[33]),
    .inData_34(stage_7_per_in[34]),
    .inData_35(stage_7_per_in[35]),
    .inData_36(stage_7_per_in[36]),
    .inData_37(stage_7_per_in[37]),
    .inData_38(stage_7_per_in[38]),
    .inData_39(stage_7_per_in[39]),
    .inData_40(stage_7_per_in[40]),
    .inData_41(stage_7_per_in[41]),
    .inData_42(stage_7_per_in[42]),
    .inData_43(stage_7_per_in[43]),
    .inData_44(stage_7_per_in[44]),
    .inData_45(stage_7_per_in[45]),
    .inData_46(stage_7_per_in[46]),
    .inData_47(stage_7_per_in[47]),
    .inData_48(stage_7_per_in[48]),
    .inData_49(stage_7_per_in[49]),
    .inData_50(stage_7_per_in[50]),
    .inData_51(stage_7_per_in[51]),
    .inData_52(stage_7_per_in[52]),
    .inData_53(stage_7_per_in[53]),
    .inData_54(stage_7_per_in[54]),
    .inData_55(stage_7_per_in[55]),
    .inData_56(stage_7_per_in[56]),
    .inData_57(stage_7_per_in[57]),
    .inData_58(stage_7_per_in[58]),
    .inData_59(stage_7_per_in[59]),
    .inData_60(stage_7_per_in[60]),
    .inData_61(stage_7_per_in[61]),
    .inData_62(stage_7_per_in[62]),
    .inData_63(stage_7_per_in[63]),
    .outData_0(stage_7_per_out[0]),
    .outData_1(stage_7_per_out[1]),
    .outData_2(stage_7_per_out[2]),
    .outData_3(stage_7_per_out[3]),
    .outData_4(stage_7_per_out[4]),
    .outData_5(stage_7_per_out[5]),
    .outData_6(stage_7_per_out[6]),
    .outData_7(stage_7_per_out[7]),
    .outData_8(stage_7_per_out[8]),
    .outData_9(stage_7_per_out[9]),
    .outData_10(stage_7_per_out[10]),
    .outData_11(stage_7_per_out[11]),
    .outData_12(stage_7_per_out[12]),
    .outData_13(stage_7_per_out[13]),
    .outData_14(stage_7_per_out[14]),
    .outData_15(stage_7_per_out[15]),
    .outData_16(stage_7_per_out[16]),
    .outData_17(stage_7_per_out[17]),
    .outData_18(stage_7_per_out[18]),
    .outData_19(stage_7_per_out[19]),
    .outData_20(stage_7_per_out[20]),
    .outData_21(stage_7_per_out[21]),
    .outData_22(stage_7_per_out[22]),
    .outData_23(stage_7_per_out[23]),
    .outData_24(stage_7_per_out[24]),
    .outData_25(stage_7_per_out[25]),
    .outData_26(stage_7_per_out[26]),
    .outData_27(stage_7_per_out[27]),
    .outData_28(stage_7_per_out[28]),
    .outData_29(stage_7_per_out[29]),
    .outData_30(stage_7_per_out[30]),
    .outData_31(stage_7_per_out[31]),
    .outData_32(stage_7_per_out[32]),
    .outData_33(stage_7_per_out[33]),
    .outData_34(stage_7_per_out[34]),
    .outData_35(stage_7_per_out[35]),
    .outData_36(stage_7_per_out[36]),
    .outData_37(stage_7_per_out[37]),
    .outData_38(stage_7_per_out[38]),
    .outData_39(stage_7_per_out[39]),
    .outData_40(stage_7_per_out[40]),
    .outData_41(stage_7_per_out[41]),
    .outData_42(stage_7_per_out[42]),
    .outData_43(stage_7_per_out[43]),
    .outData_44(stage_7_per_out[44]),
    .outData_45(stage_7_per_out[45]),
    .outData_46(stage_7_per_out[46]),
    .outData_47(stage_7_per_out[47]),
    .outData_48(stage_7_per_out[48]),
    .outData_49(stage_7_per_out[49]),
    .outData_50(stage_7_per_out[50]),
    .outData_51(stage_7_per_out[51]),
    .outData_52(stage_7_per_out[52]),
    .outData_53(stage_7_per_out[53]),
    .outData_54(stage_7_per_out[54]),
    .outData_55(stage_7_per_out[55]),
    .outData_56(stage_7_per_out[56]),
    .outData_57(stage_7_per_out[57]),
    .outData_58(stage_7_per_out[58]),
    .outData_59(stage_7_per_out[59]),
    .outData_60(stage_7_per_out[60]),
    .outData_61(stage_7_per_out[61]),
    .outData_62(stage_7_per_out[62]),
    .outData_63(stage_7_per_out[63]),
    .in_start(in_start[7]),
    .out_start(out_start[7]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 8 32 butterfly units
  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_0 (
    .x_in(stage_7_per_out[0]),
    .y_in(stage_7_per_out[1]),
    .x_out(stage_8_per_in[0]),
    .y_out(stage_8_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_1 (
    .x_in(stage_7_per_out[2]),
    .y_in(stage_7_per_out[3]),
    .x_out(stage_8_per_in[2]),
    .y_out(stage_8_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_2 (
    .x_in(stage_7_per_out[4]),
    .y_in(stage_7_per_out[5]),
    .x_out(stage_8_per_in[4]),
    .y_out(stage_8_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_3 (
    .x_in(stage_7_per_out[6]),
    .y_in(stage_7_per_out[7]),
    .x_out(stage_8_per_in[6]),
    .y_out(stage_8_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_4 (
    .x_in(stage_7_per_out[8]),
    .y_in(stage_7_per_out[9]),
    .x_out(stage_8_per_in[8]),
    .y_out(stage_8_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_5 (
    .x_in(stage_7_per_out[10]),
    .y_in(stage_7_per_out[11]),
    .x_out(stage_8_per_in[10]),
    .y_out(stage_8_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_6 (
    .x_in(stage_7_per_out[12]),
    .y_in(stage_7_per_out[13]),
    .x_out(stage_8_per_in[12]),
    .y_out(stage_8_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_7 (
    .x_in(stage_7_per_out[14]),
    .y_in(stage_7_per_out[15]),
    .x_out(stage_8_per_in[14]),
    .y_out(stage_8_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_8 (
    .x_in(stage_7_per_out[16]),
    .y_in(stage_7_per_out[17]),
    .x_out(stage_8_per_in[16]),
    .y_out(stage_8_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_9 (
    .x_in(stage_7_per_out[18]),
    .y_in(stage_7_per_out[19]),
    .x_out(stage_8_per_in[18]),
    .y_out(stage_8_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_10 (
    .x_in(stage_7_per_out[20]),
    .y_in(stage_7_per_out[21]),
    .x_out(stage_8_per_in[20]),
    .y_out(stage_8_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_11 (
    .x_in(stage_7_per_out[22]),
    .y_in(stage_7_per_out[23]),
    .x_out(stage_8_per_in[22]),
    .y_out(stage_8_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_12 (
    .x_in(stage_7_per_out[24]),
    .y_in(stage_7_per_out[25]),
    .x_out(stage_8_per_in[24]),
    .y_out(stage_8_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_13 (
    .x_in(stage_7_per_out[26]),
    .y_in(stage_7_per_out[27]),
    .x_out(stage_8_per_in[26]),
    .y_out(stage_8_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_14 (
    .x_in(stage_7_per_out[28]),
    .y_in(stage_7_per_out[29]),
    .x_out(stage_8_per_in[28]),
    .y_out(stage_8_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_15 (
    .x_in(stage_7_per_out[30]),
    .y_in(stage_7_per_out[31]),
    .x_out(stage_8_per_in[30]),
    .y_out(stage_8_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_16 (
    .x_in(stage_7_per_out[32]),
    .y_in(stage_7_per_out[33]),
    .x_out(stage_8_per_in[32]),
    .y_out(stage_8_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_17 (
    .x_in(stage_7_per_out[34]),
    .y_in(stage_7_per_out[35]),
    .x_out(stage_8_per_in[34]),
    .y_out(stage_8_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_18 (
    .x_in(stage_7_per_out[36]),
    .y_in(stage_7_per_out[37]),
    .x_out(stage_8_per_in[36]),
    .y_out(stage_8_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_19 (
    .x_in(stage_7_per_out[38]),
    .y_in(stage_7_per_out[39]),
    .x_out(stage_8_per_in[38]),
    .y_out(stage_8_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_20 (
    .x_in(stage_7_per_out[40]),
    .y_in(stage_7_per_out[41]),
    .x_out(stage_8_per_in[40]),
    .y_out(stage_8_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_21 (
    .x_in(stage_7_per_out[42]),
    .y_in(stage_7_per_out[43]),
    .x_out(stage_8_per_in[42]),
    .y_out(stage_8_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_22 (
    .x_in(stage_7_per_out[44]),
    .y_in(stage_7_per_out[45]),
    .x_out(stage_8_per_in[44]),
    .y_out(stage_8_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_23 (
    .x_in(stage_7_per_out[46]),
    .y_in(stage_7_per_out[47]),
    .x_out(stage_8_per_in[46]),
    .y_out(stage_8_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_24 (
    .x_in(stage_7_per_out[48]),
    .y_in(stage_7_per_out[49]),
    .x_out(stage_8_per_in[48]),
    .y_out(stage_8_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_25 (
    .x_in(stage_7_per_out[50]),
    .y_in(stage_7_per_out[51]),
    .x_out(stage_8_per_in[50]),
    .y_out(stage_8_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_26 (
    .x_in(stage_7_per_out[52]),
    .y_in(stage_7_per_out[53]),
    .x_out(stage_8_per_in[52]),
    .y_out(stage_8_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_27 (
    .x_in(stage_7_per_out[54]),
    .y_in(stage_7_per_out[55]),
    .x_out(stage_8_per_in[54]),
    .y_out(stage_8_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_28 (
    .x_in(stage_7_per_out[56]),
    .y_in(stage_7_per_out[57]),
    .x_out(stage_8_per_in[56]),
    .y_out(stage_8_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_29 (
    .x_in(stage_7_per_out[58]),
    .y_in(stage_7_per_out[59]),
    .x_out(stage_8_per_in[58]),
    .y_out(stage_8_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_30 (
    .x_in(stage_7_per_out[60]),
    .y_in(stage_7_per_out[61]),
    .x_out(stage_8_per_in[60]),
    .y_out(stage_8_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_31 (
    .x_in(stage_7_per_out[62]),
    .y_in(stage_7_per_out[63]),
    .x_out(stage_8_per_in[62]),
    .y_out(stage_8_per_in[63]),
    .clk(clk),
    .rst(rst)
  );



  // TODO(Yang): stage 8 -> stage 9 permutation
  // FIXME: ignore butterfly units for now.
  stage_8_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_8_9_per (
    .inData_0(stage_8_per_in[0]),
    .inData_1(stage_8_per_in[1]),
    .inData_2(stage_8_per_in[2]),
    .inData_3(stage_8_per_in[3]),
    .inData_4(stage_8_per_in[4]),
    .inData_5(stage_8_per_in[5]),
    .inData_6(stage_8_per_in[6]),
    .inData_7(stage_8_per_in[7]),
    .inData_8(stage_8_per_in[8]),
    .inData_9(stage_8_per_in[9]),
    .inData_10(stage_8_per_in[10]),
    .inData_11(stage_8_per_in[11]),
    .inData_12(stage_8_per_in[12]),
    .inData_13(stage_8_per_in[13]),
    .inData_14(stage_8_per_in[14]),
    .inData_15(stage_8_per_in[15]),
    .inData_16(stage_8_per_in[16]),
    .inData_17(stage_8_per_in[17]),
    .inData_18(stage_8_per_in[18]),
    .inData_19(stage_8_per_in[19]),
    .inData_20(stage_8_per_in[20]),
    .inData_21(stage_8_per_in[21]),
    .inData_22(stage_8_per_in[22]),
    .inData_23(stage_8_per_in[23]),
    .inData_24(stage_8_per_in[24]),
    .inData_25(stage_8_per_in[25]),
    .inData_26(stage_8_per_in[26]),
    .inData_27(stage_8_per_in[27]),
    .inData_28(stage_8_per_in[28]),
    .inData_29(stage_8_per_in[29]),
    .inData_30(stage_8_per_in[30]),
    .inData_31(stage_8_per_in[31]),
    .inData_32(stage_8_per_in[32]),
    .inData_33(stage_8_per_in[33]),
    .inData_34(stage_8_per_in[34]),
    .inData_35(stage_8_per_in[35]),
    .inData_36(stage_8_per_in[36]),
    .inData_37(stage_8_per_in[37]),
    .inData_38(stage_8_per_in[38]),
    .inData_39(stage_8_per_in[39]),
    .inData_40(stage_8_per_in[40]),
    .inData_41(stage_8_per_in[41]),
    .inData_42(stage_8_per_in[42]),
    .inData_43(stage_8_per_in[43]),
    .inData_44(stage_8_per_in[44]),
    .inData_45(stage_8_per_in[45]),
    .inData_46(stage_8_per_in[46]),
    .inData_47(stage_8_per_in[47]),
    .inData_48(stage_8_per_in[48]),
    .inData_49(stage_8_per_in[49]),
    .inData_50(stage_8_per_in[50]),
    .inData_51(stage_8_per_in[51]),
    .inData_52(stage_8_per_in[52]),
    .inData_53(stage_8_per_in[53]),
    .inData_54(stage_8_per_in[54]),
    .inData_55(stage_8_per_in[55]),
    .inData_56(stage_8_per_in[56]),
    .inData_57(stage_8_per_in[57]),
    .inData_58(stage_8_per_in[58]),
    .inData_59(stage_8_per_in[59]),
    .inData_60(stage_8_per_in[60]),
    .inData_61(stage_8_per_in[61]),
    .inData_62(stage_8_per_in[62]),
    .inData_63(stage_8_per_in[63]),
    .outData_0(stage_8_per_out[0]),
    .outData_1(stage_8_per_out[1]),
    .outData_2(stage_8_per_out[2]),
    .outData_3(stage_8_per_out[3]),
    .outData_4(stage_8_per_out[4]),
    .outData_5(stage_8_per_out[5]),
    .outData_6(stage_8_per_out[6]),
    .outData_7(stage_8_per_out[7]),
    .outData_8(stage_8_per_out[8]),
    .outData_9(stage_8_per_out[9]),
    .outData_10(stage_8_per_out[10]),
    .outData_11(stage_8_per_out[11]),
    .outData_12(stage_8_per_out[12]),
    .outData_13(stage_8_per_out[13]),
    .outData_14(stage_8_per_out[14]),
    .outData_15(stage_8_per_out[15]),
    .outData_16(stage_8_per_out[16]),
    .outData_17(stage_8_per_out[17]),
    .outData_18(stage_8_per_out[18]),
    .outData_19(stage_8_per_out[19]),
    .outData_20(stage_8_per_out[20]),
    .outData_21(stage_8_per_out[21]),
    .outData_22(stage_8_per_out[22]),
    .outData_23(stage_8_per_out[23]),
    .outData_24(stage_8_per_out[24]),
    .outData_25(stage_8_per_out[25]),
    .outData_26(stage_8_per_out[26]),
    .outData_27(stage_8_per_out[27]),
    .outData_28(stage_8_per_out[28]),
    .outData_29(stage_8_per_out[29]),
    .outData_30(stage_8_per_out[30]),
    .outData_31(stage_8_per_out[31]),
    .outData_32(stage_8_per_out[32]),
    .outData_33(stage_8_per_out[33]),
    .outData_34(stage_8_per_out[34]),
    .outData_35(stage_8_per_out[35]),
    .outData_36(stage_8_per_out[36]),
    .outData_37(stage_8_per_out[37]),
    .outData_38(stage_8_per_out[38]),
    .outData_39(stage_8_per_out[39]),
    .outData_40(stage_8_per_out[40]),
    .outData_41(stage_8_per_out[41]),
    .outData_42(stage_8_per_out[42]),
    .outData_43(stage_8_per_out[43]),
    .outData_44(stage_8_per_out[44]),
    .outData_45(stage_8_per_out[45]),
    .outData_46(stage_8_per_out[46]),
    .outData_47(stage_8_per_out[47]),
    .outData_48(stage_8_per_out[48]),
    .outData_49(stage_8_per_out[49]),
    .outData_50(stage_8_per_out[50]),
    .outData_51(stage_8_per_out[51]),
    .outData_52(stage_8_per_out[52]),
    .outData_53(stage_8_per_out[53]),
    .outData_54(stage_8_per_out[54]),
    .outData_55(stage_8_per_out[55]),
    .outData_56(stage_8_per_out[56]),
    .outData_57(stage_8_per_out[57]),
    .outData_58(stage_8_per_out[58]),
    .outData_59(stage_8_per_out[59]),
    .outData_60(stage_8_per_out[60]),
    .outData_61(stage_8_per_out[61]),
    .outData_62(stage_8_per_out[62]),
    .outData_63(stage_8_per_out[63]),
    .in_start(in_start[8]),
    .out_start(out_start[8]),
    .clk(clk),
    .rst(rst)
  );

  // TODO(Tian): stage 9 32 butterfly units
  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_0 (
    .x_in(stage_8_per_out[0]),
    .y_in(stage_8_per_out[1]),
    .x_out(stage_9_per_in[0]),
    .y_out(stage_9_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_1 (
    .x_in(stage_8_per_out[2]),
    .y_in(stage_8_per_out[3]),
    .x_out(stage_9_per_in[2]),
    .y_out(stage_9_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_2 (
    .x_in(stage_8_per_out[4]),
    .y_in(stage_8_per_out[5]),
    .x_out(stage_9_per_in[4]),
    .y_out(stage_9_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_3 (
    .x_in(stage_8_per_out[6]),
    .y_in(stage_8_per_out[7]),
    .x_out(stage_9_per_in[6]),
    .y_out(stage_9_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_4 (
    .x_in(stage_8_per_out[8]),
    .y_in(stage_8_per_out[9]),
    .x_out(stage_9_per_in[8]),
    .y_out(stage_9_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_5 (
    .x_in(stage_8_per_out[10]),
    .y_in(stage_8_per_out[11]),
    .x_out(stage_9_per_in[10]),
    .y_out(stage_9_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_6 (
    .x_in(stage_8_per_out[12]),
    .y_in(stage_8_per_out[13]),
    .x_out(stage_9_per_in[12]),
    .y_out(stage_9_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_7 (
    .x_in(stage_8_per_out[14]),
    .y_in(stage_8_per_out[15]),
    .x_out(stage_9_per_in[14]),
    .y_out(stage_9_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_8 (
    .x_in(stage_8_per_out[16]),
    .y_in(stage_8_per_out[17]),
    .x_out(stage_9_per_in[16]),
    .y_out(stage_9_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_9 (
    .x_in(stage_8_per_out[18]),
    .y_in(stage_8_per_out[19]),
    .x_out(stage_9_per_in[18]),
    .y_out(stage_9_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_10 (
    .x_in(stage_8_per_out[20]),
    .y_in(stage_8_per_out[21]),
    .x_out(stage_9_per_in[20]),
    .y_out(stage_9_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_11 (
    .x_in(stage_8_per_out[22]),
    .y_in(stage_8_per_out[23]),
    .x_out(stage_9_per_in[22]),
    .y_out(stage_9_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_12 (
    .x_in(stage_8_per_out[24]),
    .y_in(stage_8_per_out[25]),
    .x_out(stage_9_per_in[24]),
    .y_out(stage_9_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_13 (
    .x_in(stage_8_per_out[26]),
    .y_in(stage_8_per_out[27]),
    .x_out(stage_9_per_in[26]),
    .y_out(stage_9_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_14 (
    .x_in(stage_8_per_out[28]),
    .y_in(stage_8_per_out[29]),
    .x_out(stage_9_per_in[28]),
    .y_out(stage_9_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_15 (
    .x_in(stage_8_per_out[30]),
    .y_in(stage_8_per_out[31]),
    .x_out(stage_9_per_in[30]),
    .y_out(stage_9_per_in[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_16 (
    .x_in(stage_8_per_out[32]),
    .y_in(stage_8_per_out[33]),
    .x_out(stage_9_per_in[32]),
    .y_out(stage_9_per_in[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_17 (
    .x_in(stage_8_per_out[34]),
    .y_in(stage_8_per_out[35]),
    .x_out(stage_9_per_in[34]),
    .y_out(stage_9_per_in[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_18 (
    .x_in(stage_8_per_out[36]),
    .y_in(stage_8_per_out[37]),
    .x_out(stage_9_per_in[36]),
    .y_out(stage_9_per_in[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_19 (
    .x_in(stage_8_per_out[38]),
    .y_in(stage_8_per_out[39]),
    .x_out(stage_9_per_in[38]),
    .y_out(stage_9_per_in[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_20 (
    .x_in(stage_8_per_out[40]),
    .y_in(stage_8_per_out[41]),
    .x_out(stage_9_per_in[40]),
    .y_out(stage_9_per_in[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_21 (
    .x_in(stage_8_per_out[42]),
    .y_in(stage_8_per_out[43]),
    .x_out(stage_9_per_in[42]),
    .y_out(stage_9_per_in[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_22 (
    .x_in(stage_8_per_out[44]),
    .y_in(stage_8_per_out[45]),
    .x_out(stage_9_per_in[44]),
    .y_out(stage_9_per_in[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_23 (
    .x_in(stage_8_per_out[46]),
    .y_in(stage_8_per_out[47]),
    .x_out(stage_9_per_in[46]),
    .y_out(stage_9_per_in[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_24 (
    .x_in(stage_8_per_out[48]),
    .y_in(stage_8_per_out[49]),
    .x_out(stage_9_per_in[48]),
    .y_out(stage_9_per_in[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_25 (
    .x_in(stage_8_per_out[50]),
    .y_in(stage_8_per_out[51]),
    .x_out(stage_9_per_in[50]),
    .y_out(stage_9_per_in[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_26 (
    .x_in(stage_8_per_out[52]),
    .y_in(stage_8_per_out[53]),
    .x_out(stage_9_per_in[52]),
    .y_out(stage_9_per_in[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_27 (
    .x_in(stage_8_per_out[54]),
    .y_in(stage_8_per_out[55]),
    .x_out(stage_9_per_in[54]),
    .y_out(stage_9_per_in[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_28 (
    .x_in(stage_8_per_out[56]),
    .y_in(stage_8_per_out[57]),
    .x_out(stage_9_per_in[56]),
    .y_out(stage_9_per_in[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_29 (
    .x_in(stage_8_per_out[58]),
    .y_in(stage_8_per_out[59]),
    .x_out(stage_9_per_in[58]),
    .y_out(stage_9_per_in[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_30 (
    .x_in(stage_8_per_out[60]),
    .y_in(stage_8_per_out[61]),
    .x_out(stage_9_per_in[60]),
    .y_out(stage_9_per_in[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_31 (
    .x_in(stage_8_per_out[62]),
    .y_in(stage_8_per_out[63]),
    .x_out(stage_9_per_in[62]),
    .y_out(stage_9_per_in[63]),
    .clk(clk),
    .rst(rst)
  );



  // TODO(Yang): stage 8 -> stage 9 permutation
  // FIXME: ignore butterfly units for now.
  stage_9_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_9_10_per (
    .inData_0(stage_9_per_in[0]),
    .inData_1(stage_9_per_in[1]),
    .inData_2(stage_9_per_in[2]),
    .inData_3(stage_9_per_in[3]),
    .inData_4(stage_9_per_in[4]),
    .inData_5(stage_9_per_in[5]),
    .inData_6(stage_9_per_in[6]),
    .inData_7(stage_9_per_in[7]),
    .inData_8(stage_9_per_in[8]),
    .inData_9(stage_9_per_in[9]),
    .inData_10(stage_9_per_in[10]),
    .inData_11(stage_9_per_in[11]),
    .inData_12(stage_9_per_in[12]),
    .inData_13(stage_9_per_in[13]),
    .inData_14(stage_9_per_in[14]),
    .inData_15(stage_9_per_in[15]),
    .inData_16(stage_9_per_in[16]),
    .inData_17(stage_9_per_in[17]),
    .inData_18(stage_9_per_in[18]),
    .inData_19(stage_9_per_in[19]),
    .inData_20(stage_9_per_in[20]),
    .inData_21(stage_9_per_in[21]),
    .inData_22(stage_9_per_in[22]),
    .inData_23(stage_9_per_in[23]),
    .inData_24(stage_9_per_in[24]),
    .inData_25(stage_9_per_in[25]),
    .inData_26(stage_9_per_in[26]),
    .inData_27(stage_9_per_in[27]),
    .inData_28(stage_9_per_in[28]),
    .inData_29(stage_9_per_in[29]),
    .inData_30(stage_9_per_in[30]),
    .inData_31(stage_9_per_in[31]),
    .inData_32(stage_9_per_in[32]),
    .inData_33(stage_9_per_in[33]),
    .inData_34(stage_9_per_in[34]),
    .inData_35(stage_9_per_in[35]),
    .inData_36(stage_9_per_in[36]),
    .inData_37(stage_9_per_in[37]),
    .inData_38(stage_9_per_in[38]),
    .inData_39(stage_9_per_in[39]),
    .inData_40(stage_9_per_in[40]),
    .inData_41(stage_9_per_in[41]),
    .inData_42(stage_9_per_in[42]),
    .inData_43(stage_9_per_in[43]),
    .inData_44(stage_9_per_in[44]),
    .inData_45(stage_9_per_in[45]),
    .inData_46(stage_9_per_in[46]),
    .inData_47(stage_9_per_in[47]),
    .inData_48(stage_9_per_in[48]),
    .inData_49(stage_9_per_in[49]),
    .inData_50(stage_9_per_in[50]),
    .inData_51(stage_9_per_in[51]),
    .inData_52(stage_9_per_in[52]),
    .inData_53(stage_9_per_in[53]),
    .inData_54(stage_9_per_in[54]),
    .inData_55(stage_9_per_in[55]),
    .inData_56(stage_9_per_in[56]),
    .inData_57(stage_9_per_in[57]),
    .inData_58(stage_9_per_in[58]),
    .inData_59(stage_9_per_in[59]),
    .inData_60(stage_9_per_in[60]),
    .inData_61(stage_9_per_in[61]),
    .inData_62(stage_9_per_in[62]),
    .inData_63(stage_9_per_in[63]),
    .outData_0(stage_9_per_out[0]),
    .outData_1(stage_9_per_out[1]),
    .outData_2(stage_9_per_out[2]),
    .outData_3(stage_9_per_out[3]),
    .outData_4(stage_9_per_out[4]),
    .outData_5(stage_9_per_out[5]),
    .outData_6(stage_9_per_out[6]),
    .outData_7(stage_9_per_out[7]),
    .outData_8(stage_9_per_out[8]),
    .outData_9(stage_9_per_out[9]),
    .outData_10(stage_9_per_out[10]),
    .outData_11(stage_9_per_out[11]),
    .outData_12(stage_9_per_out[12]),
    .outData_13(stage_9_per_out[13]),
    .outData_14(stage_9_per_out[14]),
    .outData_15(stage_9_per_out[15]),
    .outData_16(stage_9_per_out[16]),
    .outData_17(stage_9_per_out[17]),
    .outData_18(stage_9_per_out[18]),
    .outData_19(stage_9_per_out[19]),
    .outData_20(stage_9_per_out[20]),
    .outData_21(stage_9_per_out[21]),
    .outData_22(stage_9_per_out[22]),
    .outData_23(stage_9_per_out[23]),
    .outData_24(stage_9_per_out[24]),
    .outData_25(stage_9_per_out[25]),
    .outData_26(stage_9_per_out[26]),
    .outData_27(stage_9_per_out[27]),
    .outData_28(stage_9_per_out[28]),
    .outData_29(stage_9_per_out[29]),
    .outData_30(stage_9_per_out[30]),
    .outData_31(stage_9_per_out[31]),
    .outData_32(stage_9_per_out[32]),
    .outData_33(stage_9_per_out[33]),
    .outData_34(stage_9_per_out[34]),
    .outData_35(stage_9_per_out[35]),
    .outData_36(stage_9_per_out[36]),
    .outData_37(stage_9_per_out[37]),
    .outData_38(stage_9_per_out[38]),
    .outData_39(stage_9_per_out[39]),
    .outData_40(stage_9_per_out[40]),
    .outData_41(stage_9_per_out[41]),
    .outData_42(stage_9_per_out[42]),
    .outData_43(stage_9_per_out[43]),
    .outData_44(stage_9_per_out[44]),
    .outData_45(stage_9_per_out[45]),
    .outData_46(stage_9_per_out[46]),
    .outData_47(stage_9_per_out[47]),
    .outData_48(stage_9_per_out[48]),
    .outData_49(stage_9_per_out[49]),
    .outData_50(stage_9_per_out[50]),
    .outData_51(stage_9_per_out[51]),
    .outData_52(stage_9_per_out[52]),
    .outData_53(stage_9_per_out[53]),
    .outData_54(stage_9_per_out[54]),
    .outData_55(stage_9_per_out[55]),
    .outData_56(stage_9_per_out[56]),
    .outData_57(stage_9_per_out[57]),
    .outData_58(stage_9_per_out[58]),
    .outData_59(stage_9_per_out[59]),
    .outData_60(stage_9_per_out[60]),
    .outData_61(stage_9_per_out[61]),
    .outData_62(stage_9_per_out[62]),
    .outData_63(stage_9_per_out[63]),
    .in_start(in_start[9]),
    .out_start(out_start[9]),
    .clk(clk),
    .rst(rst)
  );

  // TODO(Tian): stage 9 32 butterfly units
  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_0 (
    .x_in(stage_9_per_out[0]),
    .y_in(stage_9_per_out[1]),
    .x_out(outData[0]),
    .y_out(outData[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_1 (
    .x_in(stage_9_per_out[2]),
    .y_in(stage_9_per_out[3]),
    .x_out(outData[2]),
    .y_out(outData[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_2 (
    .x_in(stage_9_per_out[4]),
    .y_in(stage_9_per_out[5]),
    .x_out(outData[4]),
    .y_out(outData[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_3 (
    .x_in(stage_9_per_out[6]),
    .y_in(stage_9_per_out[7]),
    .x_out(outData[6]),
    .y_out(outData[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_4 (
    .x_in(stage_9_per_out[8]),
    .y_in(stage_9_per_out[9]),
    .x_out(outData[8]),
    .y_out(outData[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_5 (
    .x_in(stage_9_per_out[10]),
    .y_in(stage_9_per_out[11]),
    .x_out(outData[10]),
    .y_out(outData[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_6 (
    .x_in(stage_9_per_out[12]),
    .y_in(stage_9_per_out[13]),
    .x_out(outData[12]),
    .y_out(outData[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_7 (
    .x_in(stage_9_per_out[14]),
    .y_in(stage_9_per_out[15]),
    .x_out(outData[14]),
    .y_out(outData[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_8 (
    .x_in(stage_9_per_out[16]),
    .y_in(stage_9_per_out[17]),
    .x_out(outData[16]),
    .y_out(outData[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_9 (
    .x_in(stage_9_per_out[18]),
    .y_in(stage_9_per_out[19]),
    .x_out(outData[18]),
    .y_out(outData[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_10 (
    .x_in(stage_9_per_out[20]),
    .y_in(stage_9_per_out[21]),
    .x_out(outData[20]),
    .y_out(outData[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_11 (
    .x_in(stage_9_per_out[22]),
    .y_in(stage_9_per_out[23]),
    .x_out(outData[22]),
    .y_out(outData[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_12 (
    .x_in(stage_9_per_out[24]),
    .y_in(stage_9_per_out[25]),
    .x_out(outData[24]),
    .y_out(outData[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_13 (
    .x_in(stage_9_per_out[26]),
    .y_in(stage_9_per_out[27]),
    .x_out(outData[26]),
    .y_out(outData[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_14 (
    .x_in(stage_9_per_out[28]),
    .y_in(stage_9_per_out[29]),
    .x_out(outData[28]),
    .y_out(outData[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_15 (
    .x_in(stage_9_per_out[30]),
    .y_in(stage_9_per_out[31]),
    .x_out(outData[30]),
    .y_out(outData[31]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_16 (
    .x_in(stage_9_per_out[32]),
    .y_in(stage_9_per_out[33]),
    .x_out(outData[32]),
    .y_out(outData[33]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_17 (
    .x_in(stage_9_per_out[34]),
    .y_in(stage_9_per_out[35]),
    .x_out(outData[34]),
    .y_out(outData[35]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_18 (
    .x_in(stage_9_per_out[36]),
    .y_in(stage_9_per_out[37]),
    .x_out(outData[36]),
    .y_out(outData[37]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_19 (
    .x_in(stage_9_per_out[38]),
    .y_in(stage_9_per_out[39]),
    .x_out(outData[38]),
    .y_out(outData[39]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_20 (
    .x_in(stage_9_per_out[40]),
    .y_in(stage_9_per_out[41]),
    .x_out(outData[40]),
    .y_out(outData[41]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_21 (
    .x_in(stage_9_per_out[42]),
    .y_in(stage_9_per_out[43]),
    .x_out(outData[42]),
    .y_out(outData[43]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_22 (
    .x_in(stage_9_per_out[44]),
    .y_in(stage_9_per_out[45]),
    .x_out(outData[44]),
    .y_out(outData[45]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_23 (
    .x_in(stage_9_per_out[46]),
    .y_in(stage_9_per_out[47]),
    .x_out(outData[46]),
    .y_out(outData[47]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_24 (
    .x_in(stage_9_per_out[48]),
    .y_in(stage_9_per_out[49]),
    .x_out(outData[48]),
    .y_out(outData[49]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_25 (
    .x_in(stage_9_per_out[50]),
    .y_in(stage_9_per_out[51]),
    .x_out(outData[50]),
    .y_out(outData[51]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_26 (
    .x_in(stage_9_per_out[52]),
    .y_in(stage_9_per_out[53]),
    .x_out(outData[52]),
    .y_out(outData[53]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_27 (
    .x_in(stage_9_per_out[54]),
    .y_in(stage_9_per_out[55]),
    .x_out(outData[54]),
    .y_out(outData[55]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_28 (
    .x_in(stage_9_per_out[56]),
    .y_in(stage_9_per_out[57]),
    .x_out(outData[56]),
    .y_out(outData[57]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_29 (
    .x_in(stage_9_per_out[58]),
    .y_in(stage_9_per_out[59]),
    .x_out(outData[58]),
    .y_out(outData[59]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_30 (
    .x_in(stage_9_per_out[60]),
    .y_in(stage_9_per_out[61]),
    .x_out(outData[60]),
    .y_out(outData[61]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_31 (
    .x_in(stage_9_per_out[62]),
    .y_in(stage_9_per_out[63]),
    .x_out(outData[62]),
    .y_out(outData[63]),
    .clk(clk),
    .rst(rst)
  );


endmodule
