module stage_4_permutation #(
    parameter DATA_WIDTH_PER_INPUT = 28,
    parameter INPUT_PER_CYCLE = 64
  ) (
    inData_0,
    inData_1,
    inData_2,
    inData_3,
    inData_4,
    inData_5,
    inData_6,
    inData_7,
    inData_8,
    inData_9,
    inData_10,
    inData_11,
    inData_12,
    inData_13,
    inData_14,
    inData_15,
    inData_16,
    inData_17,
    inData_18,
    inData_19,
    inData_20,
    inData_21,
    inData_22,
    inData_23,
    inData_24,
    inData_25,
    inData_26,
    inData_27,
    inData_28,
    inData_29,
    inData_30,
    inData_31,
    inData_32,
    inData_33,
    inData_34,
    inData_35,
    inData_36,
    inData_37,
    inData_38,
    inData_39,
    inData_40,
    inData_41,
    inData_42,
    inData_43,
    inData_44,
    inData_45,
    inData_46,
    inData_47,
    inData_48,
    inData_49,
    inData_50,
    inData_51,
    inData_52,
    inData_53,
    inData_54,
    inData_55,
    inData_56,
    inData_57,
    inData_58,
    inData_59,
    inData_60,
    inData_61,
    inData_62,
    inData_63,
    inData_64,
    inData_65,
    inData_66,
    inData_67,
    inData_68,
    inData_69,
    inData_70,
    inData_71,
    inData_72,
    inData_73,
    inData_74,
    inData_75,
    inData_76,
    inData_77,
    inData_78,
    inData_79,
    inData_80,
    inData_81,
    inData_82,
    inData_83,
    inData_84,
    inData_85,
    inData_86,
    inData_87,
    inData_88,
    inData_89,
    inData_90,
    inData_91,
    inData_92,
    inData_93,
    inData_94,
    inData_95,
    inData_96,
    inData_97,
    inData_98,
    inData_99,
    inData_100,
    inData_101,
    inData_102,
    inData_103,
    inData_104,
    inData_105,
    inData_106,
    inData_107,
    inData_108,
    inData_109,
    inData_110,
    inData_111,
    inData_112,
    inData_113,
    inData_114,
    inData_115,
    inData_116,
    inData_117,
    inData_118,
    inData_119,
    inData_120,
    inData_121,
    inData_122,
    inData_123,
    inData_124,
    inData_125,
    inData_126,
    inData_127,
    outData_0,
    outData_1,
    outData_2,
    outData_3,
    outData_4,
    outData_5,
    outData_6,
    outData_7,
    outData_8,
    outData_9,
    outData_10,
    outData_11,
    outData_12,
    outData_13,
    outData_14,
    outData_15,
    outData_16,
    outData_17,
    outData_18,
    outData_19,
    outData_20,
    outData_21,
    outData_22,
    outData_23,
    outData_24,
    outData_25,
    outData_26,
    outData_27,
    outData_28,
    outData_29,
    outData_30,
    outData_31,
    outData_32,
    outData_33,
    outData_34,
    outData_35,
    outData_36,
    outData_37,
    outData_38,
    outData_39,
    outData_40,
    outData_41,
    outData_42,
    outData_43,
    outData_44,
    outData_45,
    outData_46,
    outData_47,
    outData_48,
    outData_49,
    outData_50,
    outData_51,
    outData_52,
    outData_53,
    outData_54,
    outData_55,
    outData_56,
    outData_57,
    outData_58,
    outData_59,
    outData_60,
    outData_61,
    outData_62,
    outData_63,
    outData_64,
    outData_65,
    outData_66,
    outData_67,
    outData_68,
    outData_69,
    outData_70,
    outData_71,
    outData_72,
    outData_73,
    outData_74,
    outData_75,
    outData_76,
    outData_77,
    outData_78,
    outData_79,
    outData_80,
    outData_81,
    outData_82,
    outData_83,
    outData_84,
    outData_85,
    outData_86,
    outData_87,
    outData_88,
    outData_89,
    outData_90,
    outData_91,
    outData_92,
    outData_93,
    outData_94,
    outData_95,
    outData_96,
    outData_97,
    outData_98,
    outData_99,
    outData_100,
    outData_101,
    outData_102,
    outData_103,
    outData_104,
    outData_105,
    outData_106,
    outData_107,
    outData_108,
    outData_109,
    outData_110,
    outData_111,
    outData_112,
    outData_113,
    outData_114,
    outData_115,
    outData_116,
    outData_117,
    outData_118,
    outData_119,
    outData_120,
    outData_121,
    outData_122,
    outData_123,
    outData_124,
    outData_125,
    outData_126,
    outData_127,
    in_start,
    out_start,
    clk,
    rst
  );

  input clk, rst;
  input in_start;
  output logic out_start;

  input [DATA_WIDTH_PER_INPUT-1:0] inData_0;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_1;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_2;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_3;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_4;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_5;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_6;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_7;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_8;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_9;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_10;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_11;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_12;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_13;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_14;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_15;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_16;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_17;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_18;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_19;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_20;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_21;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_22;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_23;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_24;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_25;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_26;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_27;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_28;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_29;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_30;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_31;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_32;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_33;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_34;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_35;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_36;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_37;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_38;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_39;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_40;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_41;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_42;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_43;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_44;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_45;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_46;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_47;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_48;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_49;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_50;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_51;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_52;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_53;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_54;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_55;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_56;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_57;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_58;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_59;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_60;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_61;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_62;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_63;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_64;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_65;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_66;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_67;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_68;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_69;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_70;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_71;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_72;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_73;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_74;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_75;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_76;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_77;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_78;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_79;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_80;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_81;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_82;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_83;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_84;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_85;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_86;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_87;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_88;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_89;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_90;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_91;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_92;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_93;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_94;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_95;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_96;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_97;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_98;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_99;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_100;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_101;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_102;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_103;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_104;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_105;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_106;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_107;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_108;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_109;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_110;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_111;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_112;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_113;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_114;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_115;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_116;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_117;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_118;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_119;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_120;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_121;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_122;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_123;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_124;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_125;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_126;
  input [DATA_WIDTH_PER_INPUT-1:0] inData_127;

  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_0;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_1;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_2;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_3;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_4;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_5;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_6;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_7;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_8;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_9;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_10;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_11;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_12;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_13;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_14;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_15;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_16;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_17;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_18;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_19;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_20;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_21;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_22;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_23;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_24;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_25;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_26;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_27;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_28;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_29;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_30;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_31;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_32;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_33;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_34;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_35;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_36;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_37;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_38;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_39;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_40;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_41;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_42;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_43;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_44;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_45;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_46;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_47;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_48;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_49;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_50;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_51;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_52;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_53;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_54;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_55;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_56;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_57;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_58;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_59;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_60;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_61;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_62;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_63;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_64;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_65;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_66;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_67;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_68;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_69;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_70;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_71;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_72;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_73;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_74;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_75;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_76;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_77;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_78;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_79;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_80;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_81;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_82;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_83;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_84;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_85;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_86;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_87;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_88;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_89;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_90;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_91;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_92;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_93;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_94;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_95;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_96;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_97;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_98;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_99;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_100;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_101;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_102;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_103;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_104;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_105;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_106;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_107;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_108;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_109;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_110;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_111;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_112;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_113;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_114;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_115;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_116;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_117;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_118;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_119;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_120;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_121;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_122;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_123;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_124;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_125;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_126;
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData_127;


  always_ff @ (posedge clk) begin
    if (rst) begin
      outData_0 <= 0;
      outData_1 <= 0;
      outData_2 <= 0;
      outData_3 <= 0;
      outData_4 <= 0;
      outData_5 <= 0;
      outData_6 <= 0;
      outData_7 <= 0;
      outData_8 <= 0;
      outData_9 <= 0;
      outData_10 <= 0;
      outData_11 <= 0;
      outData_12 <= 0;
      outData_13 <= 0;
      outData_14 <= 0;
      outData_15 <= 0;
      outData_16 <= 0;
      outData_17 <= 0;
      outData_18 <= 0;
      outData_19 <= 0;
      outData_20 <= 0;
      outData_21 <= 0;
      outData_22 <= 0;
      outData_23 <= 0;
      outData_24 <= 0;
      outData_25 <= 0;
      outData_26 <= 0;
      outData_27 <= 0;
      outData_28 <= 0;
      outData_29 <= 0;
      outData_30 <= 0;
      outData_31 <= 0;
      outData_32 <= 0;
      outData_33 <= 0;
      outData_34 <= 0;
      outData_35 <= 0;
      outData_36 <= 0;
      outData_37 <= 0;
      outData_38 <= 0;
      outData_39 <= 0;
      outData_40 <= 0;
      outData_41 <= 0;
      outData_42 <= 0;
      outData_43 <= 0;
      outData_44 <= 0;
      outData_45 <= 0;
      outData_46 <= 0;
      outData_47 <= 0;
      outData_48 <= 0;
      outData_49 <= 0;
      outData_50 <= 0;
      outData_51 <= 0;
      outData_52 <= 0;
      outData_53 <= 0;
      outData_54 <= 0;
      outData_55 <= 0;
      outData_56 <= 0;
      outData_57 <= 0;
      outData_58 <= 0;
      outData_59 <= 0;
      outData_60 <= 0;
      outData_61 <= 0;
      outData_62 <= 0;
      outData_63 <= 0;
      outData_64 <= 0;
      outData_65 <= 0;
      outData_66 <= 0;
      outData_67 <= 0;
      outData_68 <= 0;
      outData_69 <= 0;
      outData_70 <= 0;
      outData_71 <= 0;
      outData_72 <= 0;
      outData_73 <= 0;
      outData_74 <= 0;
      outData_75 <= 0;
      outData_76 <= 0;
      outData_77 <= 0;
      outData_78 <= 0;
      outData_79 <= 0;
      outData_80 <= 0;
      outData_81 <= 0;
      outData_82 <= 0;
      outData_83 <= 0;
      outData_84 <= 0;
      outData_85 <= 0;
      outData_86 <= 0;
      outData_87 <= 0;
      outData_88 <= 0;
      outData_89 <= 0;
      outData_90 <= 0;
      outData_91 <= 0;
      outData_92 <= 0;
      outData_93 <= 0;
      outData_94 <= 0;
      outData_95 <= 0;
      outData_96 <= 0;
      outData_97 <= 0;
      outData_98 <= 0;
      outData_99 <= 0;
      outData_100 <= 0;
      outData_101 <= 0;
      outData_102 <= 0;
      outData_103 <= 0;
      outData_104 <= 0;
      outData_105 <= 0;
      outData_106 <= 0;
      outData_107 <= 0;
      outData_108 <= 0;
      outData_109 <= 0;
      outData_110 <= 0;
      outData_111 <= 0;
      outData_112 <= 0;
      outData_113 <= 0;
      outData_114 <= 0;
      outData_115 <= 0;
      outData_116 <= 0;
      outData_117 <= 0;
      outData_118 <= 0;
      outData_119 <= 0;
      outData_120 <= 0;
      outData_121 <= 0;
      outData_122 <= 0;
      outData_123 <= 0;
      outData_124 <= 0;
      outData_125 <= 0;
      outData_126 <= 0;
      outData_127 <= 0;
    end else begin
      outData_0 <= inData_0;
      outData_1 <= inData_32;
      outData_2 <= inData_2;
      outData_3 <= inData_34;
      outData_4 <= inData_4;
      outData_5 <= inData_36;
      outData_6 <= inData_6;
      outData_7 <= inData_38;
      outData_8 <= inData_8;
      outData_9 <= inData_40;
      outData_10 <= inData_10;
      outData_11 <= inData_42;
      outData_12 <= inData_12;
      outData_13 <= inData_44;
      outData_14 <= inData_14;
      outData_15 <= inData_46;
      outData_16 <= inData_16;
      outData_17 <= inData_48;
      outData_18 <= inData_18;
      outData_19 <= inData_50;
      outData_20 <= inData_20;
      outData_21 <= inData_52;
      outData_22 <= inData_22;
      outData_23 <= inData_54;
      outData_24 <= inData_24;
      outData_25 <= inData_56;
      outData_26 <= inData_26;
      outData_27 <= inData_58;
      outData_28 <= inData_28;
      outData_29 <= inData_60;
      outData_30 <= inData_30;
      outData_31 <= inData_62;
      outData_32 <= inData_1;
      outData_33 <= inData_33;
      outData_34 <= inData_3;
      outData_35 <= inData_35;
      outData_36 <= inData_5;
      outData_37 <= inData_37;
      outData_38 <= inData_7;
      outData_39 <= inData_39;
      outData_40 <= inData_9;
      outData_41 <= inData_41;
      outData_42 <= inData_11;
      outData_43 <= inData_43;
      outData_44 <= inData_13;
      outData_45 <= inData_45;
      outData_46 <= inData_15;
      outData_47 <= inData_47;
      outData_48 <= inData_17;
      outData_49 <= inData_49;
      outData_50 <= inData_19;
      outData_51 <= inData_51;
      outData_52 <= inData_21;
      outData_53 <= inData_53;
      outData_54 <= inData_23;
      outData_55 <= inData_55;
      outData_56 <= inData_25;
      outData_57 <= inData_57;
      outData_58 <= inData_27;
      outData_59 <= inData_59;
      outData_60 <= inData_29;
      outData_61 <= inData_61;
      outData_62 <= inData_31;
      outData_63 <= inData_63;

      outData_64 <= inData_64;
      outData_65 <= inData_96;
      outData_66 <= inData_66;
      outData_67 <= inData_98;
      outData_68 <= inData_68;
      outData_69 <= inData_100;
      outData_70 <= inData_70;
      outData_71 <= inData_102;

      outData_72 <= inData_72;
      outData_73 <= inData_104;
      outData_74 <= inData_74;
      outData_75 <= inData_106;
      outData_76 <= inData_76;
      outData_77 <= inData_108;
      outData_78 <= inData_78;
      outData_79 <= inData_110;

      outData_80 <= inData_80;
      outData_81 <= inData_112;
      outData_82 <= inData_82;
      outData_83 <= inData_114;
      outData_84 <= inData_84;
      outData_85 <= inData_116;
      outData_86 <= inData_86;
      outData_87 <= inData_118;

      outData_88 <= inData_88;
      outData_89 <= inData_120;
      outData_90 <= inData_90;
      outData_91 <= inData_122;
      outData_92 <= inData_92;
      outData_93 <= inData_124;
      outData_94 <= inData_94;
      outData_95 <= inData_126;

      outData_96 <= inData_65;
      outData_97 <= inData_97;
      outData_98 <= inData_67;
      outData_99 <= inData_99;
      outData_100 <= inData_69;
      outData_101 <= inData_101;
      outData_102 <= inData_71;
      outData_103 <= inData_103;

      outData_104 <= inData_73;
      outData_105 <= inData_105;
      outData_106 <= inData_75;
      outData_107 <= inData_107;
      outData_108 <= inData_77;
      outData_109 <= inData_109;
      outData_110 <= inData_79;
      outData_111 <= inData_111;

      outData_112 <= inData_81;
      outData_113 <= inData_113;
      outData_114 <= inData_83;
      outData_115 <= inData_115;
      outData_116 <= inData_85;
      outData_117 <= inData_117;
      outData_118 <= inData_87;
      outData_119 <= inData_119;

      outData_120 <= inData_89;
      outData_121 <= inData_121;
      outData_122 <= inData_91;
      outData_123 <= inData_123;
      outData_124 <= inData_93;
      outData_125 <= inData_125;
      outData_126 <= inData_95;
      outData_127 <= inData_127;
    end
  end

endmodule
