// NTT Accelerator

module NTT_Top #(
    parameter NUM_BITS_PER_INPUT = 32
  ) (
    clk,
    rst,
    in_start,
    in_data,
    out_start,
    out_data
  );

endmodule
