// NTT Accelerator

module NTT_Top #(
    parameter DATA_WIDTH_PER_INPUT = 28,
    parameter INPUT_PER_CYCLE = 32
  ) (
    inData,
    outData,
    in_start,
    out_start,
    clk,
    rst,
  );

  input clk, rst;

  input in_start[9:0];
  output logic out_start[9:0];

  input        [DATA_WIDTH_PER_INPUT-1:0] inData[INPUT_PER_CYCLE-1:0];
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_0_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_0_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_1_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_1_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_2_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_2_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_3_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_3_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_4_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_4_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_5_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_5_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_6_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_6_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_7_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_7_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_8_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_8_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_9_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_9_per_out[INPUT_PER_CYCLE-1:0];

  parameter [7:0] START_CYCLE[11] = {0, 7, 14, 21, 28, 49, 71, 95, 123, 159, 211};

  // TODO(Tian): stage 0 32 butterfly units
  butterfly #(
    .start(START_CYCLE[0]),
    .factors({66687, 207692352, 58085086, 171518128, 153619107, 45213202, 41046131, 231691713,
              189026714, 184120139, 70631961, 79909455, 197498270, 20654843, 125081754, 22483780,
              54194127, 241662912, 186938437, 53018448, 218565763, 29126603, 176985668, 166849602,
              66993197, 242981970, 149817301, 134488788, 44349942, 215932651, 106663692, 230537579,
              209875154, 123744505, 265093046, 13110486, 243595082, 204305824, 40001367, 124635721,
              188637512, 213462715, 130849588, 188476710, 80900544, 13136617, 41376169, 134518349,
              74661667, 22903087, 9521161, 79252444, 117448591, 34884345, 216779302, 94872102,
              67400723, 110850189, 241368847, 200589425, 190155959, 7804022, 121954140, 138643341}))
  stage_0_butterfly_0 (
    .x_in(inData[0]),
    .y_in(inData[1]),
    .x_out(stage_0_per_in[0]),
    .y_out(stage_0_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({69710552, 255875272, 157049837, 60493834, 29541109, 199654780, 109238580, 264692686,
              176646986, 222469354, 66294444, 156023579, 4184358, 164354184, 261365258, 264722248,
              216344829, 224632066, 157159811, 42984958, 218464636, 10057303, 109752985, 19948338,
              107013281, 224618046, 83173794, 78067214, 82066131, 174707320, 127177690, 111544693,
              211324969, 42559975, 73580010, 58402192, 262853884, 135644103, 104968162, 29014999,
              241404981, 248367053, 127320617, 153843002, 96861137, 52859373, 111883252, 212200386,
              163120146, 114169496, 164222678, 261854403, 180135303, 98181554, 222243486, 251666562,
              47960804, 29380441, 11479903, 205236983, 185458452, 2705617, 14425613, 214088558}))
  stage_0_butterfly_1 (
    .x_in(inData[2]),
    .y_in(inData[3]),
    .x_out(stage_0_per_in[2]),
    .y_out(stage_0_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({262755833, 154212375, 25367770, 14131216, 72606471, 254000355, 131386739, 248921617,
              24152300, 43817935, 113066699, 181198907, 230614882, 168908433, 212990958, 9304145,
              83248807, 255369977, 224274217, 53103748, 56718282, 127930513, 64307891, 267667077,
              80152118, 18101390, 6554463, 152808181, 249749550, 144813234, 177333030, 120419308,
              112928859, 142863934, 103520242, 121172029, 11377467, 125480758, 212660495, 205274966,
              9977836, 177181340, 248813222, 1429580, 256522921, 153907308, 42903438, 198035948,
              243952581, 124518160, 81165688, 258225039, 13005428, 107122996, 122372515, 78535147,
              127264350, 90748831, 194452250, 48447796, 97371131, 210266721, 250007587, 25148713}))
  stage_0_butterfly_2 (
    .x_in(inData[4]),
    .y_in(inData[5]),
    .x_out(stage_0_per_in[4]),
    .y_out(stage_0_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({256317058, 5651134, 176574100, 235215540, 196552678, 65092548, 4087463, 246972075,
              197359850, 205553550, 144888817, 254205318, 116252651, 219432305, 251186267, 209423491,
              227177249, 52761187, 37869546, 77043356, 254559948, 268253695, 80396852, 243436973,
              267404879, 145663803, 243900215, 207221115, 230038199, 193252183, 186920055, 178131021,
              183986337, 153035867, 143442800, 141410653, 77239454, 209091203, 9418848, 202016934,
              136554761, 105651679, 30998042, 219873665, 234127283, 130965208, 28513237, 263341785,
              7407334, 46629005, 185511309, 119697484, 246139244, 219164507, 207114911, 200991325,
              48499686, 99140149, 132216843, 169530517, 65241583, 37489037, 13394971, 233412603}))
  stage_0_butterfly_3 (
    .x_in(inData[6]),
    .y_in(inData[7]),
    .x_out(stage_0_per_in[6]),
    .y_out(stage_0_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({36785021, 96644160, 116176624, 238066757, 241027889, 95745785, 2568552, 94477870,
              135965343, 173093264, 220939348, 20028125, 67459976, 24122396, 156421542, 145706676,
              53251080, 130184658, 139206238, 182490652, 37830528, 176845896, 85925921, 200245646,
              250343614, 75240990, 64508043, 78372181, 92664685, 175360485, 16229147, 230913482,
              259190760, 13214022, 5284602, 72907110, 178626802, 158913333, 34279912, 144340508,
              186026798, 3731063, 229577517, 193915015, 159848863, 20163279, 132170867, 143364478,
              118263349, 124384681, 183471966, 218119669, 188624074, 8903594, 35688570, 162610901,
              133533317, 224762304, 204610446, 176649880, 96783518, 101221270, 129161289, 91136142}))
  stage_0_butterfly_4 (
    .x_in(inData[8]),
    .y_in(inData[9]),
    .x_out(stage_0_per_in[8]),
    .y_out(stage_0_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({70884448, 208516738, 20380320, 156384032, 62553766, 38429557, 246330337, 18485653,
              17337072, 107466416, 259358426, 74839506, 221333762, 76096071, 79007221, 101664410,
              125436993, 155494097, 165481068, 83440545, 34758721, 24169593, 76840577, 214277734,
              119165597, 132749847, 143713813, 15448747, 57880935, 243480557, 159288788, 232016200,
              185327331, 200835165, 121708429, 150529015, 26950622, 218922070, 31628247, 176876579,
              116219557, 241656403, 64402402, 121678256, 86425411, 199114532, 210629837, 144387747,
              264754058, 75455626, 160223263, 237212534, 189299702, 56848151, 38129962, 189248627,
              112174110, 92098334, 148301509, 234435452, 75689991, 238700391, 181758089, 35697312}))
  stage_0_butterfly_5 (
    .x_in(inData[10]),
    .y_in(inData[11]),
    .x_out(stage_0_per_in[10]),
    .y_out(stage_0_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({144486207, 141475285, 33861678, 122417419, 62424622, 114175494, 171258656, 187658742,
              30978406, 41031357, 191233099, 82105625, 108814743, 76495986, 200295213, 78726832,
              240329350, 204045920, 119553807, 41015351, 17095567, 184775632, 119820987, 215044990,
              125990181, 216035935, 74620568, 100034642, 195258296, 187345691, 211474022, 123869779,
              213018760, 182322028, 217483488, 172927150, 224076531, 172413463, 124175107, 226568978,
              241147279, 81774581, 43396787, 126650083, 163686509, 64059298, 267034870, 200458300,
              21814275, 229077055, 119858575, 267701123, 233629950, 116261862, 65363597, 50041017,
              61366355, 114456140, 128923754, 28569588, 207436891, 12549924, 258398710, 113970703}))
  stage_0_butterfly_6 (
    .x_in(inData[12]),
    .y_in(inData[13]),
    .x_out(stage_0_per_in[12]),
    .y_out(stage_0_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({4869479, 250979164, 226423252, 101235253, 240913336, 219155874, 161193348, 75430495,
              7525756, 127603059, 183816509, 7373784, 45529198, 150750886, 227631635, 106279827,
              117082039, 8437385, 85943438, 241484731, 5742112, 210367757, 55952036, 50956256,
              158362238, 184194991, 114499544, 88850354, 183015243, 73886338, 224620084, 202657965,
              98446051, 222855093, 90415400, 20476611, 202037642, 117740425, 80852279, 210930243,
              219647998, 159837268, 85610695, 250769297, 35399020, 1381761, 16387901, 104273059,
              70993112, 56672741, 56349189, 15252454, 89363633, 230462114, 72373951, 260125445,
              135336752, 196403691, 211284483, 179888950, 102019874, 161018204, 212643172, 228180092}))
  stage_0_butterfly_7 (
    .x_in(inData[14]),
    .y_in(inData[15]),
    .x_out(stage_0_per_in[14]),
    .y_out(stage_0_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({181036575, 149046252, 15406607, 249303130, 118216948, 197016099, 28990836, 127667482,
              153827860, 219408463, 152434516, 90833651, 95356163, 88694916, 190584784, 154780521,
              104721465, 152028008, 207179347, 210835738, 195777196, 91129770, 62694765, 54694187,
              192617727, 233855133, 199997052, 159375180, 185375251, 89556414, 141917139, 153057061,
              171269635, 172630653, 66106013, 229787934, 236173805, 64197737, 48487396, 174554842,
              86222094, 236960516, 64123411, 144089543, 86412198, 194834330, 29149935, 182882105,
              67895486, 50484120, 111028502, 143928593, 220487343, 77305748, 129596600, 221852517,
              126869459, 60951044, 74346844, 232958416, 115863951, 185120175, 9083394, 218263368}))
  stage_0_butterfly_8 (
    .x_in(inData[16]),
    .y_in(inData[17]),
    .x_out(stage_0_per_in[16]),
    .y_out(stage_0_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({164585197, 82259521, 84197948, 196076822, 162343477, 208392312, 24580196, 205950205,
              112847505, 194382796, 104494180, 58882681, 239438610, 226909804, 195751196, 57420105,
              255042189, 104225870, 27101256, 265484036, 167135704, 162889363, 178774268, 101451720,
              126420356, 222836343, 60187882, 146642358, 92935276, 100770703, 201970932, 94729012,
              242966976, 253791818, 100723721, 11727916, 113735821, 114289273, 128081279, 122009767,
              209335538, 206932975, 55000619, 218155940, 40931981, 246263559, 3906588, 207289252,
              254651521, 50021352, 6839312, 22696094, 126673466, 74643322, 35544064, 33986901,
              257856584, 247062782, 240580313, 3059556, 218254116, 127281316, 28589493, 202839194}))
  stage_0_butterfly_9 (
    .x_in(inData[18]),
    .y_in(inData[19]),
    .x_out(stage_0_per_in[18]),
    .y_out(stage_0_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({124689641, 89494679, 12048336, 172777377, 16967674, 75161941, 165964934, 173116375,
              63479516, 209076586, 264758616, 33161823, 246348641, 52952054, 12994463, 79746145,
              151222684, 219476260, 126817458, 188253439, 15203085, 217984510, 266062977, 49412866,
              158406994, 263485445, 118812967, 263389379, 231508432, 184266218, 209775390, 116815899,
              145325214, 124256170, 115675578, 236561162, 246040827, 119485143, 131952477, 59945410,
              128639456, 214979600, 174110644, 214652925, 151896708, 218479673, 248430418, 242718809,
              43308742, 125264465, 68558047, 111988251, 186490797, 77506253, 26451456, 197145719,
              227605745, 122774092, 81924749, 130025327, 100306740, 220111512, 187430880, 80477336}))
  stage_0_butterfly_10 (
    .x_in(inData[20]),
    .y_in(inData[21]),
    .x_out(stage_0_per_in[20]),
    .y_out(stage_0_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({236609676, 108936038, 155632772, 11247416, 208367077, 12030631, 237702991, 148728622,
              192156570, 139714595, 169217935, 242696977, 111861272, 232215778, 141932586, 176645554,
              46680870, 134032627, 4080689, 253775510, 91771920, 5933624, 64186729, 204816575,
              196972136, 60114085, 24281843, 101380813, 81641436, 131659808, 120623833, 40136402,
              224193580, 41504705, 181657279, 14923017, 114906207, 1996702, 157158700, 72665107,
              66698835, 203299319, 246446391, 140980229, 15304900, 185097589, 41918325, 63912782,
              79432680, 54250256, 35256934, 172134458, 46133075, 70728737, 228992312, 37207751,
              185850221, 95857789, 34535827, 202868018, 267892175, 44186331, 94113816, 172355039}))
  stage_0_butterfly_11 (
    .x_in(inData[22]),
    .y_in(inData[23]),
    .x_out(stage_0_per_in[22]),
    .y_out(stage_0_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({175181826, 9453674, 25921170, 122635188, 129053745, 71023991, 59004276, 7487276,
              89839882, 234963902, 119598304, 99687432, 180106398, 7289546, 75588758, 195650024,
              94844905, 232700332, 232035425, 73305984, 76258087, 76831465, 194631063, 122925753,
              129973973, 136763023, 182519003, 45684920, 13646129, 170218646, 215427609, 19111856,
              111161696, 184394225, 182035415, 34093582, 143397255, 189966412, 175887545, 6456449,
              218411001, 25932042, 242432529, 207587513, 127510598, 177566022, 210485515, 148535761,
              214331009, 114664154, 124878920, 207578860, 181264550, 69161829, 103427147, 157107117,
              239446376, 14128368, 6261383, 63900610, 100616259, 126629575, 213513532, 248049881}))
  stage_0_butterfly_12 (
    .x_in(inData[24]),
    .y_in(inData[25]),
    .x_out(stage_0_per_in[24]),
    .y_out(stage_0_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({53666796, 149565630, 201841490, 229646063, 250734390, 32353046, 21867329, 94417879,
              195126393, 223749061, 18807047, 151510274, 154135831, 175735543, 96098889, 19569387,
              201750613, 179997990, 56301526, 268223107, 226796218, 176150397, 75267274, 146917464,
              215876710, 246670007, 86146205, 220989018, 242906033, 130341794, 106441080, 245173438,
              51299486, 168090046, 183906538, 133543242, 186023395, 36426289, 149121135, 32769539,
              37292607, 33343400, 66456987, 246049881, 127868408, 190924029, 95362545, 195750117,
              159083887, 83665434, 124980045, 79351768, 41512397, 71466452, 216420108, 132980811,
              35769351, 44753328, 177659362, 15241225, 254862428, 255807486, 175699854, 100791881}))
  stage_0_butterfly_13 (
    .x_in(inData[26]),
    .y_in(inData[27]),
    .x_out(stage_0_per_in[26]),
    .y_out(stage_0_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({134572374, 20490089, 54591848, 172426762, 259641163, 54291647, 266184237, 83798709,
              124903743, 240846316, 243356346, 252329804, 110349263, 106939991, 217947353, 39161232,
              260055946, 62605527, 260941520, 121709085, 39159482, 194584338, 198451374, 111058309,
              188610091, 189935724, 143647295, 177655074, 16321430, 239135625, 85861280, 121236629,
              196727396, 197999089, 4628244, 85557225, 259902883, 127312784, 176734838, 233358957,
              52172809, 222818810, 88659311, 65939487, 37689469, 35608242, 246253529, 217412044,
              263768524, 66352780, 44002169, 50385541, 153805373, 203207502, 164064761, 38583127,
              16680201, 178750844, 72006316, 178548754, 104486975, 259334239, 161494327, 85449542}))
  stage_0_butterfly_14 (
    .x_in(inData[28]),
    .y_in(inData[29]),
    .x_out(stage_0_per_in[28]),
    .y_out(stage_0_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({251547338, 198469359, 187954050, 200880844, 9599856, 107222748, 253615348, 106713399,
              145040924, 94741987, 31515852, 89730483, 75051406, 92263376, 158367942, 6208689,
              245518247, 243959994, 147907047, 132063071, 126638229, 70296940, 197375798, 91839141,
              13677670, 97932506, 208399648, 117068649, 45577615, 144316291, 102496219, 258128862,
              259597052, 244981517, 139662643, 254780782, 140652682, 75414331, 88068083, 209997049,
              22419281, 103192680, 154457559, 213843220, 209499403, 241593066, 119681087, 90431622,
              202709135, 230254857, 11713205, 92468150, 221869909, 263850390, 187446019, 231864746,
              13905102, 14195884, 61031492, 180859208, 236043136, 5071752, 81363847, 86422302}))
  stage_0_butterfly_15 (
    .x_in(inData[30]),
    .y_in(inData[31]),
    .x_out(stage_0_per_in[30]),
    .y_out(stage_0_per_in[31]),
    .clk(clk),
    .rst(rst)
  );




  // TODO(Yang): stage 0 -> stage 1 permutation
  // FIXME: ignore butterfly units for now.
  stage_0_permutation #(
    .DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    .INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_0_1_per (
    .inData_0(stage_0_per_in[0]),
    .inData_1(stage_0_per_in[1]),
    .inData_2(stage_0_per_in[2]),
    .inData_3(stage_0_per_in[3]),
    .inData_4(stage_0_per_in[4]),
    .inData_5(stage_0_per_in[5]),
    .inData_6(stage_0_per_in[6]),
    .inData_7(stage_0_per_in[7]),
    .inData_8(stage_0_per_in[8]),
    .inData_9(stage_0_per_in[9]),
    .inData_10(stage_0_per_in[10]),
    .inData_11(stage_0_per_in[11]),
    .inData_12(stage_0_per_in[12]),
    .inData_13(stage_0_per_in[13]),
    .inData_14(stage_0_per_in[14]),
    .inData_15(stage_0_per_in[15]),
    .inData_16(stage_0_per_in[16]),
    .inData_17(stage_0_per_in[17]),
    .inData_18(stage_0_per_in[18]),
    .inData_19(stage_0_per_in[19]),
    .inData_20(stage_0_per_in[20]),
    .inData_21(stage_0_per_in[21]),
    .inData_22(stage_0_per_in[22]),
    .inData_23(stage_0_per_in[23]),
    .inData_24(stage_0_per_in[24]),
    .inData_25(stage_0_per_in[25]),
    .inData_26(stage_0_per_in[26]),
    .inData_27(stage_0_per_in[27]),
    .inData_28(stage_0_per_in[28]),
    .inData_29(stage_0_per_in[29]),
    .inData_30(stage_0_per_in[30]),
    .inData_31(stage_0_per_in[31]),
    .outData_0(stage_0_per_out[0]),
    .outData_1(stage_0_per_out[1]),
    .outData_2(stage_0_per_out[2]),
    .outData_3(stage_0_per_out[3]),
    .outData_4(stage_0_per_out[4]),
    .outData_5(stage_0_per_out[5]),
    .outData_6(stage_0_per_out[6]),
    .outData_7(stage_0_per_out[7]),
    .outData_8(stage_0_per_out[8]),
    .outData_9(stage_0_per_out[9]),
    .outData_10(stage_0_per_out[10]),
    .outData_11(stage_0_per_out[11]),
    .outData_12(stage_0_per_out[12]),
    .outData_13(stage_0_per_out[13]),
    .outData_14(stage_0_per_out[14]),
    .outData_15(stage_0_per_out[15]),
    .outData_16(stage_0_per_out[16]),
    .outData_17(stage_0_per_out[17]),
    .outData_18(stage_0_per_out[18]),
    .outData_19(stage_0_per_out[19]),
    .outData_20(stage_0_per_out[20]),
    .outData_21(stage_0_per_out[21]),
    .outData_22(stage_0_per_out[22]),
    .outData_23(stage_0_per_out[23]),
    .outData_24(stage_0_per_out[24]),
    .outData_25(stage_0_per_out[25]),
    .outData_26(stage_0_per_out[26]),
    .outData_27(stage_0_per_out[27]),
    .outData_28(stage_0_per_out[28]),
    .outData_29(stage_0_per_out[29]),
    .outData_30(stage_0_per_out[30]),
    .outData_31(stage_0_per_out[31]),
    .in_start(in_start[0]),
    .out_start(out_start[0]),
    .clk(clk),
    .rst(rst)
  );

  // TODO(Tian): stage 1 32 butterfly units
  butterfly #(
    .start(START_CYCLE[1]),
    .factors({153237233, 165180840, 76624935, 99012968, 137060289, 100343421, 103368916, 29594281,
              180764097, 167181901, 265109260, 94741537, 138513718, 243339369, 232173019, 262368251,
              20917227, 146639516, 227453822, 164079161, 73099736, 84700854, 168674209, 46197346,
              44888494, 259533807, 135080569, 193174373, 121414397, 64771890, 261458154, 73072346,
              174391063, 38252193, 160856494, 81263879, 43977927, 217210388, 135902522, 102698816,
              56257750, 133952844, 172655984, 202480866, 2486257, 259164217, 82483914, 244022079,
              21253452, 108831626, 99543252, 121145061, 259302720, 23442787, 267785378, 267017218,
              128052734, 195692414, 244216061, 212728405, 205242220, 231354349, 20236367, 3021514}))
  stage_1_butterfly_0 (
    .x_in(stage_0_per_out[0]),
    .y_in(stage_0_per_out[1]),
    .x_out(stage_1_per_in[0]),
    .y_out(stage_1_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({153237233, 165180840, 76624935, 99012968, 137060289, 100343421, 103368916, 29594281,
              180764097, 167181901, 265109260, 94741537, 138513718, 243339369, 232173019, 262368251,
              20917227, 146639516, 227453822, 164079161, 73099736, 84700854, 168674209, 46197346,
              44888494, 259533807, 135080569, 193174373, 121414397, 64771890, 261458154, 73072346,
              174391063, 38252193, 160856494, 81263879, 43977927, 217210388, 135902522, 102698816,
              56257750, 133952844, 172655984, 202480866, 2486257, 259164217, 82483914, 244022079,
              21253452, 108831626, 99543252, 121145061, 259302720, 23442787, 267785378, 267017218,
              128052734, 195692414, 244216061, 212728405, 205242220, 231354349, 20236367, 3021514}))
  stage_1_butterfly_1 (
    .x_in(stage_0_per_out[2]),
    .y_in(stage_0_per_out[3]),
    .x_out(stage_1_per_in[2]),
    .y_out(stage_1_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({83809662, 168373202, 57946842, 159491687, 46312994, 73071114, 15655486, 255737752,
              172715743, 156837559, 9793208, 58491201, 160048836, 244423105, 66337349, 102243739,
              228243008, 100611174, 56207397, 1592710, 119878395, 178382895, 42575603, 189033696,
              205934027, 237395333, 59894768, 164473684, 112070980, 10310370, 159148996, 72509307,
              89028484, 54714468, 166334964, 266378632, 134161265, 98410858, 78767945, 238590283,
              21649526, 107503597, 34932582, 62027985, 112825183, 122609533, 253487730, 173513151,
              170100736, 21582278, 36492987, 107940029, 209643171, 8748458, 228572460, 7376627,
              144648965, 108164959, 232038388, 113049121, 72369588, 154317057, 171841734, 34052825}))
  stage_1_butterfly_2 (
    .x_in(stage_0_per_out[4]),
    .y_in(stage_0_per_out[5]),
    .x_out(stage_1_per_in[4]),
    .y_out(stage_1_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({83809662, 168373202, 57946842, 159491687, 46312994, 73071114, 15655486, 255737752,
              172715743, 156837559, 9793208, 58491201, 160048836, 244423105, 66337349, 102243739,
              228243008, 100611174, 56207397, 1592710, 119878395, 178382895, 42575603, 189033696,
              205934027, 237395333, 59894768, 164473684, 112070980, 10310370, 159148996, 72509307,
              89028484, 54714468, 166334964, 266378632, 134161265, 98410858, 78767945, 238590283,
              21649526, 107503597, 34932582, 62027985, 112825183, 122609533, 253487730, 173513151,
              170100736, 21582278, 36492987, 107940029, 209643171, 8748458, 228572460, 7376627,
              144648965, 108164959, 232038388, 113049121, 72369588, 154317057, 171841734, 34052825}))
  stage_1_butterfly_3 (
    .x_in(stage_0_per_out[6]),
    .y_in(stage_0_per_out[7]),
    .x_out(stage_1_per_in[6]),
    .y_out(stage_1_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({257723260, 4457103, 25278905, 121355275, 164865927, 236209279, 121608761, 79121706,
              245986816, 75689102, 85740049, 247714871, 46282885, 128011618, 82779345, 142807968,
              156534179, 259719559, 74931497, 67784869, 226025718, 169092523, 255818084, 94341361,
              76313029, 255478273, 242717180, 2204580, 249947221, 263649093, 262630184, 12817079,
              113006603, 50606491, 175949223, 122969043, 187381670, 202871094, 188535281, 248922055,
              234775081, 214937778, 90701762, 207877484, 217359458, 201160126, 94178347, 149904904,
              248946430, 110378476, 267860193, 70033082, 191242693, 195152646, 44896056, 104557844,
              10943590, 86359417, 136898494, 39337018, 87202745, 240930884, 237616434, 128159746}))
  stage_1_butterfly_4 (
    .x_in(stage_0_per_out[8]),
    .y_in(stage_0_per_out[9]),
    .x_out(stage_1_per_in[8]),
    .y_out(stage_1_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({257723260, 4457103, 25278905, 121355275, 164865927, 236209279, 121608761, 79121706,
              245986816, 75689102, 85740049, 247714871, 46282885, 128011618, 82779345, 142807968,
              156534179, 259719559, 74931497, 67784869, 226025718, 169092523, 255818084, 94341361,
              76313029, 255478273, 242717180, 2204580, 249947221, 263649093, 262630184, 12817079,
              113006603, 50606491, 175949223, 122969043, 187381670, 202871094, 188535281, 248922055,
              234775081, 214937778, 90701762, 207877484, 217359458, 201160126, 94178347, 149904904,
              248946430, 110378476, 267860193, 70033082, 191242693, 195152646, 44896056, 104557844,
              10943590, 86359417, 136898494, 39337018, 87202745, 240930884, 237616434, 128159746}))
  stage_1_butterfly_5 (
    .x_in(stage_0_per_out[10]),
    .y_in(stage_0_per_out[11]),
    .x_out(stage_1_per_in[10]),
    .y_out(stage_1_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({267008435, 248328138, 65803974, 112174557, 198352904, 12711531, 133573372, 230871518,
              53126225, 254234203, 211646222, 128995628, 185175266, 161607031, 233083676, 118444917,
              207021189, 218195682, 219133933, 148649408, 78273516, 217993137, 67241659, 148479452,
              138629310, 82321748, 143811089, 24036023, 13228372, 187988754, 122025398, 132747224,
              18793692, 184464011, 155613159, 173577844, 45457492, 1807449, 116513948, 120217110,
              99899421, 86350556, 31964447, 118320134, 198957507, 188526794, 116527240, 184177651,
              53025186, 115050087, 232740066, 186476418, 146205579, 207530748, 50523873, 7226699,
              264322432, 1855205, 16351380, 7280660, 159987098, 189909138, 165584204, 123018041}))
  stage_1_butterfly_6 (
    .x_in(stage_0_per_out[12]),
    .y_in(stage_0_per_out[13]),
    .x_out(stage_1_per_in[12]),
    .y_out(stage_1_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({267008435, 248328138, 65803974, 112174557, 198352904, 12711531, 133573372, 230871518,
              53126225, 254234203, 211646222, 128995628, 185175266, 161607031, 233083676, 118444917,
              207021189, 218195682, 219133933, 148649408, 78273516, 217993137, 67241659, 148479452,
              138629310, 82321748, 143811089, 24036023, 13228372, 187988754, 122025398, 132747224,
              18793692, 184464011, 155613159, 173577844, 45457492, 1807449, 116513948, 120217110,
              99899421, 86350556, 31964447, 118320134, 198957507, 188526794, 116527240, 184177651,
              53025186, 115050087, 232740066, 186476418, 146205579, 207530748, 50523873, 7226699,
              264322432, 1855205, 16351380, 7280660, 159987098, 189909138, 165584204, 123018041}))
  stage_1_butterfly_7 (
    .x_in(stage_0_per_out[14]),
    .y_in(stage_0_per_out[15]),
    .x_out(stage_1_per_in[14]),
    .y_out(stage_1_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({181617487, 207769332, 5445105, 36213609, 167645260, 34402629, 266777383, 136179523,
              215525211, 120466187, 210373784, 184522009, 69017626, 246741831, 193451294, 135921552,
              243047656, 62094530, 211824237, 259895089, 5267255, 234786570, 206844979, 64464693,
              18433789, 127918992, 40915578, 100027171, 12912005, 263648524, 139742686, 241071152,
              83977288, 248251528, 125713617, 133098101, 62456195, 73481957, 251672258, 198043993,
              127163336, 81414740, 74458128, 209744644, 175710456, 187208958, 230865684, 190453366,
              176911171, 30998914, 151857114, 32319537, 146399832, 263725948, 169792793, 54916848,
              44047649, 245372433, 45355620, 128297265, 205604517, 110720332, 129677075, 23586243}))
  stage_1_butterfly_8 (
    .x_in(stage_0_per_out[16]),
    .y_in(stage_0_per_out[17]),
    .x_out(stage_1_per_in[16]),
    .y_out(stage_1_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({181617487, 207769332, 5445105, 36213609, 167645260, 34402629, 266777383, 136179523,
              215525211, 120466187, 210373784, 184522009, 69017626, 246741831, 193451294, 135921552,
              243047656, 62094530, 211824237, 259895089, 5267255, 234786570, 206844979, 64464693,
              18433789, 127918992, 40915578, 100027171, 12912005, 263648524, 139742686, 241071152,
              83977288, 248251528, 125713617, 133098101, 62456195, 73481957, 251672258, 198043993,
              127163336, 81414740, 74458128, 209744644, 175710456, 187208958, 230865684, 190453366,
              176911171, 30998914, 151857114, 32319537, 146399832, 263725948, 169792793, 54916848,
              44047649, 245372433, 45355620, 128297265, 205604517, 110720332, 129677075, 23586243}))
  stage_1_butterfly_9 (
    .x_in(stage_0_per_out[18]),
    .y_in(stage_0_per_out[19]),
    .x_out(stage_1_per_in[18]),
    .y_out(stage_1_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({3395282, 164728317, 36620312, 115053845, 77119896, 110055875, 195181845, 145831337,
              249311139, 204707946, 87492030, 101783683, 108319109, 212788230, 129694458, 218380292,
              19700796, 209780385, 62513408, 54393228, 199055975, 92902456, 215085706, 174856430,
              7301415, 19817676, 11850588, 98445813, 116257755, 141267184, 133565368, 209154967,
              194684542, 222249559, 157839041, 144502563, 64830196, 84669572, 17682401, 139101859,
              43819650, 104121890, 236272786, 121712648, 12286825, 26068775, 182803613, 104215821,
              94436408, 2487567, 238832783, 216819035, 84798700, 105443909, 226834391, 97171493,
              209708523, 134561032, 70944317, 138215130, 141562255, 120261431, 133273987, 248732744}))
  stage_1_butterfly_10 (
    .x_in(stage_0_per_out[20]),
    .y_in(stage_0_per_out[21]),
    .x_out(stage_1_per_in[20]),
    .y_out(stage_1_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({3395282, 164728317, 36620312, 115053845, 77119896, 110055875, 195181845, 145831337,
              249311139, 204707946, 87492030, 101783683, 108319109, 212788230, 129694458, 218380292,
              19700796, 209780385, 62513408, 54393228, 199055975, 92902456, 215085706, 174856430,
              7301415, 19817676, 11850588, 98445813, 116257755, 141267184, 133565368, 209154967,
              194684542, 222249559, 157839041, 144502563, 64830196, 84669572, 17682401, 139101859,
              43819650, 104121890, 236272786, 121712648, 12286825, 26068775, 182803613, 104215821,
              94436408, 2487567, 238832783, 216819035, 84798700, 105443909, 226834391, 97171493,
              209708523, 134561032, 70944317, 138215130, 141562255, 120261431, 133273987, 248732744}))
  stage_1_butterfly_11 (
    .x_in(stage_0_per_out[22]),
    .y_in(stage_0_per_out[23]),
    .x_out(stage_1_per_in[22]),
    .y_out(stage_1_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({66412546, 206116619, 17758040, 151297332, 69205492, 128589211, 105793954, 45842328,
              224922683, 268043824, 98139687, 236829199, 244004517, 236528116, 40741603, 17642100,
              213678985, 58671364, 226759664, 183613005, 91397014, 107152911, 94686133, 55222727,
              74472522, 158067861, 112360014, 113269084, 47531240, 145317914, 203850982, 37377133,
              60051251, 18205961, 50162577, 212287973, 219484262, 33096679, 232847226, 102230592,
              16652121, 189044804, 196018390, 23328014, 56132215, 863665, 90149574, 209112367,
              50083600, 148051010, 154298223, 256834872, 106743034, 211201491, 139044757, 93757293,
              149788353, 187172755, 97163404, 159978713, 265496406, 158914825, 77783793, 263207998}))
  stage_1_butterfly_12 (
    .x_in(stage_0_per_out[24]),
    .y_in(stage_0_per_out[25]),
    .x_out(stage_1_per_in[24]),
    .y_out(stage_1_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({66412546, 206116619, 17758040, 151297332, 69205492, 128589211, 105793954, 45842328,
              224922683, 268043824, 98139687, 236829199, 244004517, 236528116, 40741603, 17642100,
              213678985, 58671364, 226759664, 183613005, 91397014, 107152911, 94686133, 55222727,
              74472522, 158067861, 112360014, 113269084, 47531240, 145317914, 203850982, 37377133,
              60051251, 18205961, 50162577, 212287973, 219484262, 33096679, 232847226, 102230592,
              16652121, 189044804, 196018390, 23328014, 56132215, 863665, 90149574, 209112367,
              50083600, 148051010, 154298223, 256834872, 106743034, 211201491, 139044757, 93757293,
              149788353, 187172755, 97163404, 159978713, 265496406, 158914825, 77783793, 263207998}))
  stage_1_butterfly_13 (
    .x_in(stage_0_per_out[26]),
    .y_in(stage_0_per_out[27]),
    .x_out(stage_1_per_in[26]),
    .y_out(stage_1_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({3341663, 207047180, 157386503, 126749676, 190540901, 142941966, 229954056, 187867192,
              90687088, 123335487, 226981541, 183590673, 211982342, 174290656, 175990762, 31243956,
              18338102, 23776027, 260110386, 94206887, 107024087, 92770973, 81838336, 12591284,
              136710753, 122455193, 255463943, 118946466, 263001722, 189816962, 101579460, 212425161,
              163823140, 163197321, 160539079, 107138937, 2017030, 77536776, 86776671, 62688241,
              228715598, 58903295, 25360705, 6257752, 126413069, 197065781, 19904170, 6828726,
              77804235, 201787732, 120080647, 43000087, 238468357, 10967191, 92441360, 75993973,
              78612624, 145056180, 254842567, 6760936, 172401093, 51838504, 79230237, 55947412}))
  stage_1_butterfly_14 (
    .x_in(stage_0_per_out[28]),
    .y_in(stage_0_per_out[29]),
    .x_out(stage_1_per_in[28]),
    .y_out(stage_1_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({3341663, 207047180, 157386503, 126749676, 190540901, 142941966, 229954056, 187867192,
              90687088, 123335487, 226981541, 183590673, 211982342, 174290656, 175990762, 31243956,
              18338102, 23776027, 260110386, 94206887, 107024087, 92770973, 81838336, 12591284,
              136710753, 122455193, 255463943, 118946466, 263001722, 189816962, 101579460, 212425161,
              163823140, 163197321, 160539079, 107138937, 2017030, 77536776, 86776671, 62688241,
              228715598, 58903295, 25360705, 6257752, 126413069, 197065781, 19904170, 6828726,
              77804235, 201787732, 120080647, 43000087, 238468357, 10967191, 92441360, 75993973,
              78612624, 145056180, 254842567, 6760936, 172401093, 51838504, 79230237, 55947412}))
  stage_1_butterfly_15 (
    .x_in(stage_0_per_out[30]),
    .y_in(stage_0_per_out[31]),
    .x_out(stage_1_per_in[30]),
    .y_out(stage_1_per_in[31]),
    .clk(clk),
    .rst(rst)
  );




  
  // TODO(Yang): stage 1 -> stage 2 permutation
  // FIXME: ignore butterfly units for now.
  stage_1_permutation #(
    .DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    .INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_1_2_per (
    .inData_0(stage_1_per_in[0]),
    .inData_1(stage_1_per_in[1]),
    .inData_2(stage_1_per_in[2]),
    .inData_3(stage_1_per_in[3]),
    .inData_4(stage_1_per_in[4]),
    .inData_5(stage_1_per_in[5]),
    .inData_6(stage_1_per_in[6]),
    .inData_7(stage_1_per_in[7]),
    .inData_8(stage_1_per_in[8]),
    .inData_9(stage_1_per_in[9]),
    .inData_10(stage_1_per_in[10]),
    .inData_11(stage_1_per_in[11]),
    .inData_12(stage_1_per_in[12]),
    .inData_13(stage_1_per_in[13]),
    .inData_14(stage_1_per_in[14]),
    .inData_15(stage_1_per_in[15]),
    .inData_16(stage_1_per_in[16]),
    .inData_17(stage_1_per_in[17]),
    .inData_18(stage_1_per_in[18]),
    .inData_19(stage_1_per_in[19]),
    .inData_20(stage_1_per_in[20]),
    .inData_21(stage_1_per_in[21]),
    .inData_22(stage_1_per_in[22]),
    .inData_23(stage_1_per_in[23]),
    .inData_24(stage_1_per_in[24]),
    .inData_25(stage_1_per_in[25]),
    .inData_26(stage_1_per_in[26]),
    .inData_27(stage_1_per_in[27]),
    .inData_28(stage_1_per_in[28]),
    .inData_29(stage_1_per_in[29]),
    .inData_30(stage_1_per_in[30]),
    .inData_31(stage_1_per_in[31]),
    .outData_0(stage_1_per_out[0]),
    .outData_1(stage_1_per_out[1]),
    .outData_2(stage_1_per_out[2]),
    .outData_3(stage_1_per_out[3]),
    .outData_4(stage_1_per_out[4]),
    .outData_5(stage_1_per_out[5]),
    .outData_6(stage_1_per_out[6]),
    .outData_7(stage_1_per_out[7]),
    .outData_8(stage_1_per_out[8]),
    .outData_9(stage_1_per_out[9]),
    .outData_10(stage_1_per_out[10]),
    .outData_11(stage_1_per_out[11]),
    .outData_12(stage_1_per_out[12]),
    .outData_13(stage_1_per_out[13]),
    .outData_14(stage_1_per_out[14]),
    .outData_15(stage_1_per_out[15]),
    .outData_16(stage_1_per_out[16]),
    .outData_17(stage_1_per_out[17]),
    .outData_18(stage_1_per_out[18]),
    .outData_19(stage_1_per_out[19]),
    .outData_20(stage_1_per_out[20]),
    .outData_21(stage_1_per_out[21]),
    .outData_22(stage_1_per_out[22]),
    .outData_23(stage_1_per_out[23]),
    .outData_24(stage_1_per_out[24]),
    .outData_25(stage_1_per_out[25]),
    .outData_26(stage_1_per_out[26]),
    .outData_27(stage_1_per_out[27]),
    .outData_28(stage_1_per_out[28]),
    .outData_29(stage_1_per_out[29]),
    .outData_30(stage_1_per_out[30]),
    .outData_31(stage_1_per_out[31]),
    .in_start(in_start[1]),
    .out_start(out_start[1]),
    .clk(clk),
    .rst(rst)
  );


  // TODO(Tian): stage 2 32 butterfly units
  butterfly #(
    .start(START_CYCLE[2]),
    .factors({184644727, 21080194, 171051327, 126063290, 43104106, 145034471, 224225395, 256272276,
              196522490, 44547301, 167366585, 219083512, 218147185, 166955734, 213835479, 237102043,
              193915204, 218231468, 165350229, 175719113, 206705681, 61997323, 117507527, 156366160,
              242516310, 49504466, 158168844, 36946189, 165872957, 11500489, 261795000, 95861179,
              98085790, 169480001, 67225153, 202071175, 42355602, 34481514, 28242170, 222683851,
              186863562, 136992892, 259958064, 225650462, 109479656, 205961920, 182702557, 62844488,
              242425786, 187864761, 131304314, 266671862, 82155735, 95282463, 55609416, 59284831,
              141424302, 5292226, 118377542, 95560742, 92160417, 136878682, 56246211, 138879618}))
  stage_2_butterfly_0 (
    .x_in(stage_1_per_out[0]),
    .y_in(stage_1_per_out[1]),
    .x_out(stage_2_per_in[0]),
    .y_out(stage_2_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({184644727, 21080194, 171051327, 126063290, 43104106, 145034471, 224225395, 256272276,
              196522490, 44547301, 167366585, 219083512, 218147185, 166955734, 213835479, 237102043,
              193915204, 218231468, 165350229, 175719113, 206705681, 61997323, 117507527, 156366160,
              242516310, 49504466, 158168844, 36946189, 165872957, 11500489, 261795000, 95861179,
              98085790, 169480001, 67225153, 202071175, 42355602, 34481514, 28242170, 222683851,
              186863562, 136992892, 259958064, 225650462, 109479656, 205961920, 182702557, 62844488,
              242425786, 187864761, 131304314, 266671862, 82155735, 95282463, 55609416, 59284831,
              141424302, 5292226, 118377542, 95560742, 92160417, 136878682, 56246211, 138879618}))
  stage_2_butterfly_1 (
    .x_in(stage_1_per_out[2]),
    .y_in(stage_1_per_out[3]),
    .x_out(stage_2_per_in[2]),
    .y_out(stage_2_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({184644727, 21080194, 171051327, 126063290, 43104106, 145034471, 224225395, 256272276,
              196522490, 44547301, 167366585, 219083512, 218147185, 166955734, 213835479, 237102043,
              193915204, 218231468, 165350229, 175719113, 206705681, 61997323, 117507527, 156366160,
              242516310, 49504466, 158168844, 36946189, 165872957, 11500489, 261795000, 95861179,
              98085790, 169480001, 67225153, 202071175, 42355602, 34481514, 28242170, 222683851,
              186863562, 136992892, 259958064, 225650462, 109479656, 205961920, 182702557, 62844488,
              242425786, 187864761, 131304314, 266671862, 82155735, 95282463, 55609416, 59284831,
              141424302, 5292226, 118377542, 95560742, 92160417, 136878682, 56246211, 138879618}))
  stage_2_butterfly_2 (
    .x_in(stage_1_per_out[4]),
    .y_in(stage_1_per_out[5]),
    .x_out(stage_2_per_in[4]),
    .y_out(stage_2_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({184644727, 21080194, 171051327, 126063290, 43104106, 145034471, 224225395, 256272276,
              196522490, 44547301, 167366585, 219083512, 218147185, 166955734, 213835479, 237102043,
              193915204, 218231468, 165350229, 175719113, 206705681, 61997323, 117507527, 156366160,
              242516310, 49504466, 158168844, 36946189, 165872957, 11500489, 261795000, 95861179,
              98085790, 169480001, 67225153, 202071175, 42355602, 34481514, 28242170, 222683851,
              186863562, 136992892, 259958064, 225650462, 109479656, 205961920, 182702557, 62844488,
              242425786, 187864761, 131304314, 266671862, 82155735, 95282463, 55609416, 59284831,
              141424302, 5292226, 118377542, 95560742, 92160417, 136878682, 56246211, 138879618}))
  stage_2_butterfly_3 (
    .x_in(stage_1_per_out[6]),
    .y_in(stage_1_per_out[7]),
    .x_out(stage_2_per_in[6]),
    .y_out(stage_2_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({255286072, 220490426, 173118058, 97439895, 185138250, 93740850, 134269022, 146037274,
              222861227, 58483920, 200399539, 206649748, 82684352, 219898221, 69584498, 10720790,
              87202272, 251138298, 29987725, 210914061, 21739535, 200749611, 171362072, 143779572,
              119169851, 73698550, 215146927, 262077011, 244477824, 242025902, 26067051, 234350511,
              135886841, 78649100, 160841949, 216395023, 135618975, 263530653, 157966005, 126520315,
              210795202, 79136411, 14568946, 224586596, 82934386, 193296437, 100123291, 191444307,
              251384491, 207329882, 40550456, 243024363, 262464837, 212214167, 217383280, 144929841,
              206252403, 58644800, 199810586, 148390399, 129576773, 209658551, 32087335, 206725018}))
  stage_2_butterfly_4 (
    .x_in(stage_1_per_out[8]),
    .y_in(stage_1_per_out[9]),
    .x_out(stage_2_per_in[8]),
    .y_out(stage_2_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({255286072, 220490426, 173118058, 97439895, 185138250, 93740850, 134269022, 146037274,
              222861227, 58483920, 200399539, 206649748, 82684352, 219898221, 69584498, 10720790,
              87202272, 251138298, 29987725, 210914061, 21739535, 200749611, 171362072, 143779572,
              119169851, 73698550, 215146927, 262077011, 244477824, 242025902, 26067051, 234350511,
              135886841, 78649100, 160841949, 216395023, 135618975, 263530653, 157966005, 126520315,
              210795202, 79136411, 14568946, 224586596, 82934386, 193296437, 100123291, 191444307,
              251384491, 207329882, 40550456, 243024363, 262464837, 212214167, 217383280, 144929841,
              206252403, 58644800, 199810586, 148390399, 129576773, 209658551, 32087335, 206725018}))
  stage_2_butterfly_5 (
    .x_in(stage_1_per_out[10]),
    .y_in(stage_1_per_out[11]),
    .x_out(stage_2_per_in[10]),
    .y_out(stage_2_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({255286072, 220490426, 173118058, 97439895, 185138250, 93740850, 134269022, 146037274,
              222861227, 58483920, 200399539, 206649748, 82684352, 219898221, 69584498, 10720790,
              87202272, 251138298, 29987725, 210914061, 21739535, 200749611, 171362072, 143779572,
              119169851, 73698550, 215146927, 262077011, 244477824, 242025902, 26067051, 234350511,
              135886841, 78649100, 160841949, 216395023, 135618975, 263530653, 157966005, 126520315,
              210795202, 79136411, 14568946, 224586596, 82934386, 193296437, 100123291, 191444307,
              251384491, 207329882, 40550456, 243024363, 262464837, 212214167, 217383280, 144929841,
              206252403, 58644800, 199810586, 148390399, 129576773, 209658551, 32087335, 206725018}))
  stage_2_butterfly_6 (
    .x_in(stage_1_per_out[12]),
    .y_in(stage_1_per_out[13]),
    .x_out(stage_2_per_in[12]),
    .y_out(stage_2_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({255286072, 220490426, 173118058, 97439895, 185138250, 93740850, 134269022, 146037274,
              222861227, 58483920, 200399539, 206649748, 82684352, 219898221, 69584498, 10720790,
              87202272, 251138298, 29987725, 210914061, 21739535, 200749611, 171362072, 143779572,
              119169851, 73698550, 215146927, 262077011, 244477824, 242025902, 26067051, 234350511,
              135886841, 78649100, 160841949, 216395023, 135618975, 263530653, 157966005, 126520315,
              210795202, 79136411, 14568946, 224586596, 82934386, 193296437, 100123291, 191444307,
              251384491, 207329882, 40550456, 243024363, 262464837, 212214167, 217383280, 144929841,
              206252403, 58644800, 199810586, 148390399, 129576773, 209658551, 32087335, 206725018}))
  stage_2_butterfly_7 (
    .x_in(stage_1_per_out[14]),
    .y_in(stage_1_per_out[15]),
    .x_out(stage_2_per_in[14]),
    .y_out(stage_2_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({158466952, 225389748, 196328787, 164638888, 34971158, 9810331, 81527994, 165134943,
              174900371, 74093574, 32260862, 18298478, 249146534, 137346680, 233514072, 10143115,
              47375162, 154421517, 124400051, 8950678, 161171966, 232451599, 202776751, 225175773,
              218694662, 43078133, 201863951, 182691070, 158727274, 247253507, 209583375, 42156432,
              102915173, 126188511, 134877507, 100457939, 169508713, 24688427, 23405380, 12196542,
              100229847, 168676526, 160254284, 234113027, 63079505, 44301230, 244763177, 65413984,
              40158424, 84058929, 181468172, 113309038, 77389872, 10003248, 219312182, 69773246,
              9842125, 68267735, 67321994, 85252512, 207821787, 188517169, 262540431, 140366124}))
  stage_2_butterfly_8 (
    .x_in(stage_1_per_out[16]),
    .y_in(stage_1_per_out[17]),
    .x_out(stage_2_per_in[16]),
    .y_out(stage_2_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({158466952, 225389748, 196328787, 164638888, 34971158, 9810331, 81527994, 165134943,
              174900371, 74093574, 32260862, 18298478, 249146534, 137346680, 233514072, 10143115,
              47375162, 154421517, 124400051, 8950678, 161171966, 232451599, 202776751, 225175773,
              218694662, 43078133, 201863951, 182691070, 158727274, 247253507, 209583375, 42156432,
              102915173, 126188511, 134877507, 100457939, 169508713, 24688427, 23405380, 12196542,
              100229847, 168676526, 160254284, 234113027, 63079505, 44301230, 244763177, 65413984,
              40158424, 84058929, 181468172, 113309038, 77389872, 10003248, 219312182, 69773246,
              9842125, 68267735, 67321994, 85252512, 207821787, 188517169, 262540431, 140366124}))
  stage_2_butterfly_9 (
    .x_in(stage_1_per_out[18]),
    .y_in(stage_1_per_out[19]),
    .x_out(stage_2_per_in[18]),
    .y_out(stage_2_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({158466952, 225389748, 196328787, 164638888, 34971158, 9810331, 81527994, 165134943,
              174900371, 74093574, 32260862, 18298478, 249146534, 137346680, 233514072, 10143115,
              47375162, 154421517, 124400051, 8950678, 161171966, 232451599, 202776751, 225175773,
              218694662, 43078133, 201863951, 182691070, 158727274, 247253507, 209583375, 42156432,
              102915173, 126188511, 134877507, 100457939, 169508713, 24688427, 23405380, 12196542,
              100229847, 168676526, 160254284, 234113027, 63079505, 44301230, 244763177, 65413984,
              40158424, 84058929, 181468172, 113309038, 77389872, 10003248, 219312182, 69773246,
              9842125, 68267735, 67321994, 85252512, 207821787, 188517169, 262540431, 140366124}))
  stage_2_butterfly_10 (
    .x_in(stage_1_per_out[20]),
    .y_in(stage_1_per_out[21]),
    .x_out(stage_2_per_in[20]),
    .y_out(stage_2_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({158466952, 225389748, 196328787, 164638888, 34971158, 9810331, 81527994, 165134943,
              174900371, 74093574, 32260862, 18298478, 249146534, 137346680, 233514072, 10143115,
              47375162, 154421517, 124400051, 8950678, 161171966, 232451599, 202776751, 225175773,
              218694662, 43078133, 201863951, 182691070, 158727274, 247253507, 209583375, 42156432,
              102915173, 126188511, 134877507, 100457939, 169508713, 24688427, 23405380, 12196542,
              100229847, 168676526, 160254284, 234113027, 63079505, 44301230, 244763177, 65413984,
              40158424, 84058929, 181468172, 113309038, 77389872, 10003248, 219312182, 69773246,
              9842125, 68267735, 67321994, 85252512, 207821787, 188517169, 262540431, 140366124}))
  stage_2_butterfly_11 (
    .x_in(stage_1_per_out[22]),
    .y_in(stage_1_per_out[23]),
    .x_out(stage_2_per_in[22]),
    .y_out(stage_2_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({160807241, 206795535, 177340471, 10112777, 199876762, 16471674, 125267062, 63483304,
              260909397, 64764693, 229100654, 172935357, 1562592, 57599709, 55567611, 66310724,
              43575145, 40718170, 252241817, 176665584, 237438985, 56943278, 42585458, 171541778,
              129101436, 244216783, 60072008, 257269778, 1613379, 232445568, 130696933, 262358962,
              99187435, 35754446, 250508912, 254132077, 77981460, 219738759, 178386996, 68736878,
              181295312, 87088032, 64884498, 5299132, 56094099, 117221766, 13458851, 190319963,
              20857483, 72621624, 27056737, 85340443, 114486793, 94612904, 196771169, 65324949,
              61345534, 57635675, 66242139, 119568150, 151095818, 192832423, 168977833, 73081523}))
  stage_2_butterfly_12 (
    .x_in(stage_1_per_out[24]),
    .y_in(stage_1_per_out[25]),
    .x_out(stage_2_per_in[24]),
    .y_out(stage_2_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({160807241, 206795535, 177340471, 10112777, 199876762, 16471674, 125267062, 63483304,
              260909397, 64764693, 229100654, 172935357, 1562592, 57599709, 55567611, 66310724,
              43575145, 40718170, 252241817, 176665584, 237438985, 56943278, 42585458, 171541778,
              129101436, 244216783, 60072008, 257269778, 1613379, 232445568, 130696933, 262358962,
              99187435, 35754446, 250508912, 254132077, 77981460, 219738759, 178386996, 68736878,
              181295312, 87088032, 64884498, 5299132, 56094099, 117221766, 13458851, 190319963,
              20857483, 72621624, 27056737, 85340443, 114486793, 94612904, 196771169, 65324949,
              61345534, 57635675, 66242139, 119568150, 151095818, 192832423, 168977833, 73081523}))
  stage_2_butterfly_13 (
    .x_in(stage_1_per_out[26]),
    .y_in(stage_1_per_out[27]),
    .x_out(stage_2_per_in[26]),
    .y_out(stage_2_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({160807241, 206795535, 177340471, 10112777, 199876762, 16471674, 125267062, 63483304,
              260909397, 64764693, 229100654, 172935357, 1562592, 57599709, 55567611, 66310724,
              43575145, 40718170, 252241817, 176665584, 237438985, 56943278, 42585458, 171541778,
              129101436, 244216783, 60072008, 257269778, 1613379, 232445568, 130696933, 262358962,
              99187435, 35754446, 250508912, 254132077, 77981460, 219738759, 178386996, 68736878,
              181295312, 87088032, 64884498, 5299132, 56094099, 117221766, 13458851, 190319963,
              20857483, 72621624, 27056737, 85340443, 114486793, 94612904, 196771169, 65324949,
              61345534, 57635675, 66242139, 119568150, 151095818, 192832423, 168977833, 73081523}))
  stage_2_butterfly_14 (
    .x_in(stage_1_per_out[28]),
    .y_in(stage_1_per_out[29]),
    .x_out(stage_2_per_in[28]),
    .y_out(stage_2_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({160807241, 206795535, 177340471, 10112777, 199876762, 16471674, 125267062, 63483304,
              260909397, 64764693, 229100654, 172935357, 1562592, 57599709, 55567611, 66310724,
              43575145, 40718170, 252241817, 176665584, 237438985, 56943278, 42585458, 171541778,
              129101436, 244216783, 60072008, 257269778, 1613379, 232445568, 130696933, 262358962,
              99187435, 35754446, 250508912, 254132077, 77981460, 219738759, 178386996, 68736878,
              181295312, 87088032, 64884498, 5299132, 56094099, 117221766, 13458851, 190319963,
              20857483, 72621624, 27056737, 85340443, 114486793, 94612904, 196771169, 65324949,
              61345534, 57635675, 66242139, 119568150, 151095818, 192832423, 168977833, 73081523}))
  stage_2_butterfly_15 (
    .x_in(stage_1_per_out[30]),
    .y_in(stage_1_per_out[31]),
    .x_out(stage_2_per_in[30]),
    .y_out(stage_2_per_in[31]),
    .clk(clk),
    .rst(rst)
  );





  // TODO(Yang): stage 2 -> stage 3 permutation
  // FIXME: ignore butterfly units for now.
  stage_2_permutation #(
    .DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    .INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_2_3_per (
    .inData_0(stage_2_per_in[0]),
    .inData_1(stage_2_per_in[1]),
    .inData_2(stage_2_per_in[2]),
    .inData_3(stage_2_per_in[3]),
    .inData_4(stage_2_per_in[4]),
    .inData_5(stage_2_per_in[5]),
    .inData_6(stage_2_per_in[6]),
    .inData_7(stage_2_per_in[7]),
    .inData_8(stage_2_per_in[8]),
    .inData_9(stage_2_per_in[9]),
    .inData_10(stage_2_per_in[10]),
    .inData_11(stage_2_per_in[11]),
    .inData_12(stage_2_per_in[12]),
    .inData_13(stage_2_per_in[13]),
    .inData_14(stage_2_per_in[14]),
    .inData_15(stage_2_per_in[15]),
    .inData_16(stage_2_per_in[16]),
    .inData_17(stage_2_per_in[17]),
    .inData_18(stage_2_per_in[18]),
    .inData_19(stage_2_per_in[19]),
    .inData_20(stage_2_per_in[20]),
    .inData_21(stage_2_per_in[21]),
    .inData_22(stage_2_per_in[22]),
    .inData_23(stage_2_per_in[23]),
    .inData_24(stage_2_per_in[24]),
    .inData_25(stage_2_per_in[25]),
    .inData_26(stage_2_per_in[26]),
    .inData_27(stage_2_per_in[27]),
    .inData_28(stage_2_per_in[28]),
    .inData_29(stage_2_per_in[29]),
    .inData_30(stage_2_per_in[30]),
    .inData_31(stage_2_per_in[31]),
    .outData_0(stage_2_per_out[0]),
    .outData_1(stage_2_per_out[1]),
    .outData_2(stage_2_per_out[2]),
    .outData_3(stage_2_per_out[3]),
    .outData_4(stage_2_per_out[4]),
    .outData_5(stage_2_per_out[5]),
    .outData_6(stage_2_per_out[6]),
    .outData_7(stage_2_per_out[7]),
    .outData_8(stage_2_per_out[8]),
    .outData_9(stage_2_per_out[9]),
    .outData_10(stage_2_per_out[10]),
    .outData_11(stage_2_per_out[11]),
    .outData_12(stage_2_per_out[12]),
    .outData_13(stage_2_per_out[13]),
    .outData_14(stage_2_per_out[14]),
    .outData_15(stage_2_per_out[15]),
    .outData_16(stage_2_per_out[16]),
    .outData_17(stage_2_per_out[17]),
    .outData_18(stage_2_per_out[18]),
    .outData_19(stage_2_per_out[19]),
    .outData_20(stage_2_per_out[20]),
    .outData_21(stage_2_per_out[21]),
    .outData_22(stage_2_per_out[22]),
    .outData_23(stage_2_per_out[23]),
    .outData_24(stage_2_per_out[24]),
    .outData_25(stage_2_per_out[25]),
    .outData_26(stage_2_per_out[26]),
    .outData_27(stage_2_per_out[27]),
    .outData_28(stage_2_per_out[28]),
    .outData_29(stage_2_per_out[29]),
    .outData_30(stage_2_per_out[30]),
    .outData_31(stage_2_per_out[31]),
    .in_start(in_start[2]),
    .out_start(out_start[2]),
    .clk(clk),
    .rst(rst)
  );

  // TODO(Tian): stage 3 32 butterfly units
  butterfly #(
    .start(START_CYCLE[3]),
    .factors({163812837, 149528048, 41086336, 163585105, 77337691, 201357873, 246744565, 161827885,
              44942358, 108810259, 63703579, 40553702, 202221416, 229216409, 212648666, 252952333,
              242800442, 211668928, 210298252, 147433882, 99962405, 248876054, 13519489, 15927889,
              98878775, 28824907, 96648403, 217644581, 184226747, 230702770, 22541719, 69161747,
              186413553, 189762285, 7055647, 133081916, 188210893, 249640399, 71064168, 257268473,
              101839787, 240677074, 119707826, 216143425, 170604387, 123185272, 257798138, 227894900,
              78777967, 63350037, 59208162, 37936257, 91898237, 241125460, 139182289, 81777479,
              183348420, 34339674, 9757140, 173702965, 250166212, 150873005, 108965460, 130557622}))
  stage_3_butterfly_0 (
    .x_in(stage_2_per_out[0]),
    .y_in(stage_2_per_out[1]),
    .x_out(stage_3_per_in[0]),
    .y_out(stage_3_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({163812837, 149528048, 41086336, 163585105, 77337691, 201357873, 246744565, 161827885,
              44942358, 108810259, 63703579, 40553702, 202221416, 229216409, 212648666, 252952333,
              242800442, 211668928, 210298252, 147433882, 99962405, 248876054, 13519489, 15927889,
              98878775, 28824907, 96648403, 217644581, 184226747, 230702770, 22541719, 69161747,
              186413553, 189762285, 7055647, 133081916, 188210893, 249640399, 71064168, 257268473,
              101839787, 240677074, 119707826, 216143425, 170604387, 123185272, 257798138, 227894900,
              78777967, 63350037, 59208162, 37936257, 91898237, 241125460, 139182289, 81777479,
              183348420, 34339674, 9757140, 173702965, 250166212, 150873005, 108965460, 130557622}))
  stage_3_butterfly_1 (
    .x_in(stage_2_per_out[2]),
    .y_in(stage_2_per_out[3]),
    .x_out(stage_3_per_in[2]),
    .y_out(stage_3_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({163812837, 149528048, 41086336, 163585105, 77337691, 201357873, 246744565, 161827885,
              44942358, 108810259, 63703579, 40553702, 202221416, 229216409, 212648666, 252952333,
              242800442, 211668928, 210298252, 147433882, 99962405, 248876054, 13519489, 15927889,
              98878775, 28824907, 96648403, 217644581, 184226747, 230702770, 22541719, 69161747,
              186413553, 189762285, 7055647, 133081916, 188210893, 249640399, 71064168, 257268473,
              101839787, 240677074, 119707826, 216143425, 170604387, 123185272, 257798138, 227894900,
              78777967, 63350037, 59208162, 37936257, 91898237, 241125460, 139182289, 81777479,
              183348420, 34339674, 9757140, 173702965, 250166212, 150873005, 108965460, 130557622}))
  stage_3_butterfly_2 (
    .x_in(stage_2_per_out[4]),
    .y_in(stage_2_per_out[5]),
    .x_out(stage_3_per_in[4]),
    .y_out(stage_3_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({163812837, 149528048, 41086336, 163585105, 77337691, 201357873, 246744565, 161827885,
              44942358, 108810259, 63703579, 40553702, 202221416, 229216409, 212648666, 252952333,
              242800442, 211668928, 210298252, 147433882, 99962405, 248876054, 13519489, 15927889,
              98878775, 28824907, 96648403, 217644581, 184226747, 230702770, 22541719, 69161747,
              186413553, 189762285, 7055647, 133081916, 188210893, 249640399, 71064168, 257268473,
              101839787, 240677074, 119707826, 216143425, 170604387, 123185272, 257798138, 227894900,
              78777967, 63350037, 59208162, 37936257, 91898237, 241125460, 139182289, 81777479,
              183348420, 34339674, 9757140, 173702965, 250166212, 150873005, 108965460, 130557622}))
  stage_3_butterfly_3 (
    .x_in(stage_2_per_out[6]),
    .y_in(stage_2_per_out[7]),
    .x_out(stage_3_per_in[6]),
    .y_out(stage_3_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({163812837, 149528048, 41086336, 163585105, 77337691, 201357873, 246744565, 161827885,
              44942358, 108810259, 63703579, 40553702, 202221416, 229216409, 212648666, 252952333,
              242800442, 211668928, 210298252, 147433882, 99962405, 248876054, 13519489, 15927889,
              98878775, 28824907, 96648403, 217644581, 184226747, 230702770, 22541719, 69161747,
              186413553, 189762285, 7055647, 133081916, 188210893, 249640399, 71064168, 257268473,
              101839787, 240677074, 119707826, 216143425, 170604387, 123185272, 257798138, 227894900,
              78777967, 63350037, 59208162, 37936257, 91898237, 241125460, 139182289, 81777479,
              183348420, 34339674, 9757140, 173702965, 250166212, 150873005, 108965460, 130557622}))
  stage_3_butterfly_4 (
    .x_in(stage_2_per_out[8]),
    .y_in(stage_2_per_out[9]),
    .x_out(stage_3_per_in[8]),
    .y_out(stage_3_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({163812837, 149528048, 41086336, 163585105, 77337691, 201357873, 246744565, 161827885,
              44942358, 108810259, 63703579, 40553702, 202221416, 229216409, 212648666, 252952333,
              242800442, 211668928, 210298252, 147433882, 99962405, 248876054, 13519489, 15927889,
              98878775, 28824907, 96648403, 217644581, 184226747, 230702770, 22541719, 69161747,
              186413553, 189762285, 7055647, 133081916, 188210893, 249640399, 71064168, 257268473,
              101839787, 240677074, 119707826, 216143425, 170604387, 123185272, 257798138, 227894900,
              78777967, 63350037, 59208162, 37936257, 91898237, 241125460, 139182289, 81777479,
              183348420, 34339674, 9757140, 173702965, 250166212, 150873005, 108965460, 130557622}))
  stage_3_butterfly_5 (
    .x_in(stage_2_per_out[10]),
    .y_in(stage_2_per_out[11]),
    .x_out(stage_3_per_in[10]),
    .y_out(stage_3_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({163812837, 149528048, 41086336, 163585105, 77337691, 201357873, 246744565, 161827885,
              44942358, 108810259, 63703579, 40553702, 202221416, 229216409, 212648666, 252952333,
              242800442, 211668928, 210298252, 147433882, 99962405, 248876054, 13519489, 15927889,
              98878775, 28824907, 96648403, 217644581, 184226747, 230702770, 22541719, 69161747,
              186413553, 189762285, 7055647, 133081916, 188210893, 249640399, 71064168, 257268473,
              101839787, 240677074, 119707826, 216143425, 170604387, 123185272, 257798138, 227894900,
              78777967, 63350037, 59208162, 37936257, 91898237, 241125460, 139182289, 81777479,
              183348420, 34339674, 9757140, 173702965, 250166212, 150873005, 108965460, 130557622}))
  stage_3_butterfly_6 (
    .x_in(stage_2_per_out[12]),
    .y_in(stage_2_per_out[13]),
    .x_out(stage_3_per_in[12]),
    .y_out(stage_3_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({163812837, 149528048, 41086336, 163585105, 77337691, 201357873, 246744565, 161827885,
              44942358, 108810259, 63703579, 40553702, 202221416, 229216409, 212648666, 252952333,
              242800442, 211668928, 210298252, 147433882, 99962405, 248876054, 13519489, 15927889,
              98878775, 28824907, 96648403, 217644581, 184226747, 230702770, 22541719, 69161747,
              186413553, 189762285, 7055647, 133081916, 188210893, 249640399, 71064168, 257268473,
              101839787, 240677074, 119707826, 216143425, 170604387, 123185272, 257798138, 227894900,
              78777967, 63350037, 59208162, 37936257, 91898237, 241125460, 139182289, 81777479,
              183348420, 34339674, 9757140, 173702965, 250166212, 150873005, 108965460, 130557622}))
  stage_3_butterfly_7 (
    .x_in(stage_2_per_out[14]),
    .y_in(stage_2_per_out[15]),
    .x_out(stage_3_per_in[14]),
    .y_out(stage_3_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({155168409, 172227818, 133503098, 3883583, 34119889, 41630462, 164195239, 2795054,
              234890903, 214551729, 241682233, 149851545, 204152715, 160286792, 254509489, 220618744,
              146361539, 144414946, 197074908, 42733001, 132703565, 258649698, 47994339, 162031725,
              258923154, 139555205, 195631434, 18399308, 196436059, 143969713, 13250338, 87844233,
              176917280, 246656426, 244883276, 238498066, 261793746, 151968102, 101483624, 68136911,
              12328961, 265950570, 39141691, 86730411, 13919506, 85922744, 170227406, 253827407,
              22463657, 214085592, 236144340, 37011073, 83853696, 25065602, 10130658, 78488715,
              106640438, 41155851, 59283803, 90597117, 100484142, 193371292, 75673633, 231318087}))
  stage_3_butterfly_8 (
    .x_in(stage_2_per_out[16]),
    .y_in(stage_2_per_out[17]),
    .x_out(stage_3_per_in[16]),
    .y_out(stage_3_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({155168409, 172227818, 133503098, 3883583, 34119889, 41630462, 164195239, 2795054,
              234890903, 214551729, 241682233, 149851545, 204152715, 160286792, 254509489, 220618744,
              146361539, 144414946, 197074908, 42733001, 132703565, 258649698, 47994339, 162031725,
              258923154, 139555205, 195631434, 18399308, 196436059, 143969713, 13250338, 87844233,
              176917280, 246656426, 244883276, 238498066, 261793746, 151968102, 101483624, 68136911,
              12328961, 265950570, 39141691, 86730411, 13919506, 85922744, 170227406, 253827407,
              22463657, 214085592, 236144340, 37011073, 83853696, 25065602, 10130658, 78488715,
              106640438, 41155851, 59283803, 90597117, 100484142, 193371292, 75673633, 231318087}))
  stage_3_butterfly_9 (
    .x_in(stage_2_per_out[18]),
    .y_in(stage_2_per_out[19]),
    .x_out(stage_3_per_in[18]),
    .y_out(stage_3_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({155168409, 172227818, 133503098, 3883583, 34119889, 41630462, 164195239, 2795054,
              234890903, 214551729, 241682233, 149851545, 204152715, 160286792, 254509489, 220618744,
              146361539, 144414946, 197074908, 42733001, 132703565, 258649698, 47994339, 162031725,
              258923154, 139555205, 195631434, 18399308, 196436059, 143969713, 13250338, 87844233,
              176917280, 246656426, 244883276, 238498066, 261793746, 151968102, 101483624, 68136911,
              12328961, 265950570, 39141691, 86730411, 13919506, 85922744, 170227406, 253827407,
              22463657, 214085592, 236144340, 37011073, 83853696, 25065602, 10130658, 78488715,
              106640438, 41155851, 59283803, 90597117, 100484142, 193371292, 75673633, 231318087}))
  stage_3_butterfly_10 (
    .x_in(stage_2_per_out[20]),
    .y_in(stage_2_per_out[21]),
    .x_out(stage_3_per_in[20]),
    .y_out(stage_3_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({155168409, 172227818, 133503098, 3883583, 34119889, 41630462, 164195239, 2795054,
              234890903, 214551729, 241682233, 149851545, 204152715, 160286792, 254509489, 220618744,
              146361539, 144414946, 197074908, 42733001, 132703565, 258649698, 47994339, 162031725,
              258923154, 139555205, 195631434, 18399308, 196436059, 143969713, 13250338, 87844233,
              176917280, 246656426, 244883276, 238498066, 261793746, 151968102, 101483624, 68136911,
              12328961, 265950570, 39141691, 86730411, 13919506, 85922744, 170227406, 253827407,
              22463657, 214085592, 236144340, 37011073, 83853696, 25065602, 10130658, 78488715,
              106640438, 41155851, 59283803, 90597117, 100484142, 193371292, 75673633, 231318087}))
  stage_3_butterfly_11 (
    .x_in(stage_2_per_out[22]),
    .y_in(stage_2_per_out[23]),
    .x_out(stage_3_per_in[22]),
    .y_out(stage_3_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({155168409, 172227818, 133503098, 3883583, 34119889, 41630462, 164195239, 2795054,
              234890903, 214551729, 241682233, 149851545, 204152715, 160286792, 254509489, 220618744,
              146361539, 144414946, 197074908, 42733001, 132703565, 258649698, 47994339, 162031725,
              258923154, 139555205, 195631434, 18399308, 196436059, 143969713, 13250338, 87844233,
              176917280, 246656426, 244883276, 238498066, 261793746, 151968102, 101483624, 68136911,
              12328961, 265950570, 39141691, 86730411, 13919506, 85922744, 170227406, 253827407,
              22463657, 214085592, 236144340, 37011073, 83853696, 25065602, 10130658, 78488715,
              106640438, 41155851, 59283803, 90597117, 100484142, 193371292, 75673633, 231318087}))
  stage_3_butterfly_12 (
    .x_in(stage_2_per_out[24]),
    .y_in(stage_2_per_out[25]),
    .x_out(stage_3_per_in[24]),
    .y_out(stage_3_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({155168409, 172227818, 133503098, 3883583, 34119889, 41630462, 164195239, 2795054,
              234890903, 214551729, 241682233, 149851545, 204152715, 160286792, 254509489, 220618744,
              146361539, 144414946, 197074908, 42733001, 132703565, 258649698, 47994339, 162031725,
              258923154, 139555205, 195631434, 18399308, 196436059, 143969713, 13250338, 87844233,
              176917280, 246656426, 244883276, 238498066, 261793746, 151968102, 101483624, 68136911,
              12328961, 265950570, 39141691, 86730411, 13919506, 85922744, 170227406, 253827407,
              22463657, 214085592, 236144340, 37011073, 83853696, 25065602, 10130658, 78488715,
              106640438, 41155851, 59283803, 90597117, 100484142, 193371292, 75673633, 231318087}))
  stage_3_butterfly_13 (
    .x_in(stage_2_per_out[26]),
    .y_in(stage_2_per_out[27]),
    .x_out(stage_3_per_in[26]),
    .y_out(stage_3_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({155168409, 172227818, 133503098, 3883583, 34119889, 41630462, 164195239, 2795054,
              234890903, 214551729, 241682233, 149851545, 204152715, 160286792, 254509489, 220618744,
              146361539, 144414946, 197074908, 42733001, 132703565, 258649698, 47994339, 162031725,
              258923154, 139555205, 195631434, 18399308, 196436059, 143969713, 13250338, 87844233,
              176917280, 246656426, 244883276, 238498066, 261793746, 151968102, 101483624, 68136911,
              12328961, 265950570, 39141691, 86730411, 13919506, 85922744, 170227406, 253827407,
              22463657, 214085592, 236144340, 37011073, 83853696, 25065602, 10130658, 78488715,
              106640438, 41155851, 59283803, 90597117, 100484142, 193371292, 75673633, 231318087}))
  stage_3_butterfly_14 (
    .x_in(stage_2_per_out[28]),
    .y_in(stage_2_per_out[29]),
    .x_out(stage_3_per_in[28]),
    .y_out(stage_3_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({155168409, 172227818, 133503098, 3883583, 34119889, 41630462, 164195239, 2795054,
              234890903, 214551729, 241682233, 149851545, 204152715, 160286792, 254509489, 220618744,
              146361539, 144414946, 197074908, 42733001, 132703565, 258649698, 47994339, 162031725,
              258923154, 139555205, 195631434, 18399308, 196436059, 143969713, 13250338, 87844233,
              176917280, 246656426, 244883276, 238498066, 261793746, 151968102, 101483624, 68136911,
              12328961, 265950570, 39141691, 86730411, 13919506, 85922744, 170227406, 253827407,
              22463657, 214085592, 236144340, 37011073, 83853696, 25065602, 10130658, 78488715,
              106640438, 41155851, 59283803, 90597117, 100484142, 193371292, 75673633, 231318087}))
  stage_3_butterfly_15 (
    .x_in(stage_2_per_out[30]),
    .y_in(stage_2_per_out[31]),
    .x_out(stage_3_per_in[30]),
    .y_out(stage_3_per_in[31]),
    .clk(clk),
    .rst(rst)
  );





  // TODO(Yang): stage 3 -> stage 4 permutation
  // FIXME: ignore butterfly units for now.
  stage_3_permutation #(
    .DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    .INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_3_4_per (
    .inData_0(stage_3_per_in[0]),
    .inData_1(stage_3_per_in[1]),
    .inData_2(stage_3_per_in[2]),
    .inData_3(stage_3_per_in[3]),
    .inData_4(stage_3_per_in[4]),
    .inData_5(stage_3_per_in[5]),
    .inData_6(stage_3_per_in[6]),
    .inData_7(stage_3_per_in[7]),
    .inData_8(stage_3_per_in[8]),
    .inData_9(stage_3_per_in[9]),
    .inData_10(stage_3_per_in[10]),
    .inData_11(stage_3_per_in[11]),
    .inData_12(stage_3_per_in[12]),
    .inData_13(stage_3_per_in[13]),
    .inData_14(stage_3_per_in[14]),
    .inData_15(stage_3_per_in[15]),
    .inData_16(stage_3_per_in[16]),
    .inData_17(stage_3_per_in[17]),
    .inData_18(stage_3_per_in[18]),
    .inData_19(stage_3_per_in[19]),
    .inData_20(stage_3_per_in[20]),
    .inData_21(stage_3_per_in[21]),
    .inData_22(stage_3_per_in[22]),
    .inData_23(stage_3_per_in[23]),
    .inData_24(stage_3_per_in[24]),
    .inData_25(stage_3_per_in[25]),
    .inData_26(stage_3_per_in[26]),
    .inData_27(stage_3_per_in[27]),
    .inData_28(stage_3_per_in[28]),
    .inData_29(stage_3_per_in[29]),
    .inData_30(stage_3_per_in[30]),
    .inData_31(stage_3_per_in[31]),
    .outData_0(stage_3_per_out[0]),
    .outData_1(stage_3_per_out[1]),
    .outData_2(stage_3_per_out[2]),
    .outData_3(stage_3_per_out[3]),
    .outData_4(stage_3_per_out[4]),
    .outData_5(stage_3_per_out[5]),
    .outData_6(stage_3_per_out[6]),
    .outData_7(stage_3_per_out[7]),
    .outData_8(stage_3_per_out[8]),
    .outData_9(stage_3_per_out[9]),
    .outData_10(stage_3_per_out[10]),
    .outData_11(stage_3_per_out[11]),
    .outData_12(stage_3_per_out[12]),
    .outData_13(stage_3_per_out[13]),
    .outData_14(stage_3_per_out[14]),
    .outData_15(stage_3_per_out[15]),
    .outData_16(stage_3_per_out[16]),
    .outData_17(stage_3_per_out[17]),
    .outData_18(stage_3_per_out[18]),
    .outData_19(stage_3_per_out[19]),
    .outData_20(stage_3_per_out[20]),
    .outData_21(stage_3_per_out[21]),
    .outData_22(stage_3_per_out[22]),
    .outData_23(stage_3_per_out[23]),
    .outData_24(stage_3_per_out[24]),
    .outData_25(stage_3_per_out[25]),
    .outData_26(stage_3_per_out[26]),
    .outData_27(stage_3_per_out[27]),
    .outData_28(stage_3_per_out[28]),
    .outData_29(stage_3_per_out[29]),
    .outData_30(stage_3_per_out[30]),
    .outData_31(stage_3_per_out[31]),
    .in_start(in_start[3]),
    .out_start(out_start[3]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 4 32 butterfly units
  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 197787791, 215696667, 172642311, 153962078, 11695616, 233560477, 189907315,
              181852808, 147699054, 146694818, 202366126, 218546733, 78852289, 227611463, 71460019,
              17079898, 193045667, 25574347, 66112528, 263678998, 115957373, 27685019, 47317233,
              179817683, 109553202, 6323336, 165226744, 200054106, 191662816, 170752771, 140204941,
              141548072, 169276669, 70982951, 119224607, 124918999, 82771912, 39593842, 239095400,
              102065274, 157085730, 109254766, 208403048, 237620966, 111341228, 210568560, 177255039,
              76642651, 41084242, 201062854, 130295133, 152865265, 175609590, 62045777, 118939950,
              168270865, 71471012, 235204060, 131798756, 162373432, 74680748, 112472991, 145384235}))
  stage_4_butterfly_0 (
    .x_in(stage_3_per_out[0]),
    .y_in(stage_3_per_out[1]),
    .x_out(stage_4_per_in[0]),
    .y_out(stage_4_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 197787791, 215696667, 172642311, 153962078, 11695616, 233560477, 189907315,
              181852808, 147699054, 146694818, 202366126, 218546733, 78852289, 227611463, 71460019,
              17079898, 193045667, 25574347, 66112528, 263678998, 115957373, 27685019, 47317233,
              179817683, 109553202, 6323336, 165226744, 200054106, 191662816, 170752771, 140204941,
              141548072, 169276669, 70982951, 119224607, 124918999, 82771912, 39593842, 239095400,
              102065274, 157085730, 109254766, 208403048, 237620966, 111341228, 210568560, 177255039,
              76642651, 41084242, 201062854, 130295133, 152865265, 175609590, 62045777, 118939950,
              168270865, 71471012, 235204060, 131798756, 162373432, 74680748, 112472991, 145384235}))
  stage_4_butterfly_1 (
    .x_in(stage_3_per_out[2]),
    .y_in(stage_3_per_out[3]),
    .x_out(stage_4_per_in[2]),
    .y_out(stage_4_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 197787791, 215696667, 172642311, 153962078, 11695616, 233560477, 189907315,
              181852808, 147699054, 146694818, 202366126, 218546733, 78852289, 227611463, 71460019,
              17079898, 193045667, 25574347, 66112528, 263678998, 115957373, 27685019, 47317233,
              179817683, 109553202, 6323336, 165226744, 200054106, 191662816, 170752771, 140204941,
              141548072, 169276669, 70982951, 119224607, 124918999, 82771912, 39593842, 239095400,
              102065274, 157085730, 109254766, 208403048, 237620966, 111341228, 210568560, 177255039,
              76642651, 41084242, 201062854, 130295133, 152865265, 175609590, 62045777, 118939950,
              168270865, 71471012, 235204060, 131798756, 162373432, 74680748, 112472991, 145384235}))
  stage_4_butterfly_2 (
    .x_in(stage_3_per_out[4]),
    .y_in(stage_3_per_out[5]),
    .x_out(stage_4_per_in[4]),
    .y_out(stage_4_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 197787791, 215696667, 172642311, 153962078, 11695616, 233560477, 189907315,
              181852808, 147699054, 146694818, 202366126, 218546733, 78852289, 227611463, 71460019,
              17079898, 193045667, 25574347, 66112528, 263678998, 115957373, 27685019, 47317233,
              179817683, 109553202, 6323336, 165226744, 200054106, 191662816, 170752771, 140204941,
              141548072, 169276669, 70982951, 119224607, 124918999, 82771912, 39593842, 239095400,
              102065274, 157085730, 109254766, 208403048, 237620966, 111341228, 210568560, 177255039,
              76642651, 41084242, 201062854, 130295133, 152865265, 175609590, 62045777, 118939950,
              168270865, 71471012, 235204060, 131798756, 162373432, 74680748, 112472991, 145384235}))
  stage_4_butterfly_3 (
    .x_in(stage_3_per_out[6]),
    .y_in(stage_3_per_out[7]),
    .x_out(stage_4_per_in[6]),
    .y_out(stage_4_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 197787791, 215696667, 172642311, 153962078, 11695616, 233560477, 189907315,
              181852808, 147699054, 146694818, 202366126, 218546733, 78852289, 227611463, 71460019,
              17079898, 193045667, 25574347, 66112528, 263678998, 115957373, 27685019, 47317233,
              179817683, 109553202, 6323336, 165226744, 200054106, 191662816, 170752771, 140204941,
              141548072, 169276669, 70982951, 119224607, 124918999, 82771912, 39593842, 239095400,
              102065274, 157085730, 109254766, 208403048, 237620966, 111341228, 210568560, 177255039,
              76642651, 41084242, 201062854, 130295133, 152865265, 175609590, 62045777, 118939950,
              168270865, 71471012, 235204060, 131798756, 162373432, 74680748, 112472991, 145384235}))
  stage_4_butterfly_4 (
    .x_in(stage_3_per_out[8]),
    .y_in(stage_3_per_out[9]),
    .x_out(stage_4_per_in[8]),
    .y_out(stage_4_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 197787791, 215696667, 172642311, 153962078, 11695616, 233560477, 189907315,
              181852808, 147699054, 146694818, 202366126, 218546733, 78852289, 227611463, 71460019,
              17079898, 193045667, 25574347, 66112528, 263678998, 115957373, 27685019, 47317233,
              179817683, 109553202, 6323336, 165226744, 200054106, 191662816, 170752771, 140204941,
              141548072, 169276669, 70982951, 119224607, 124918999, 82771912, 39593842, 239095400,
              102065274, 157085730, 109254766, 208403048, 237620966, 111341228, 210568560, 177255039,
              76642651, 41084242, 201062854, 130295133, 152865265, 175609590, 62045777, 118939950,
              168270865, 71471012, 235204060, 131798756, 162373432, 74680748, 112472991, 145384235}))
  stage_4_butterfly_5 (
    .x_in(stage_3_per_out[10]),
    .y_in(stage_3_per_out[11]),
    .x_out(stage_4_per_in[10]),
    .y_out(stage_4_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 197787791, 215696667, 172642311, 153962078, 11695616, 233560477, 189907315,
              181852808, 147699054, 146694818, 202366126, 218546733, 78852289, 227611463, 71460019,
              17079898, 193045667, 25574347, 66112528, 263678998, 115957373, 27685019, 47317233,
              179817683, 109553202, 6323336, 165226744, 200054106, 191662816, 170752771, 140204941,
              141548072, 169276669, 70982951, 119224607, 124918999, 82771912, 39593842, 239095400,
              102065274, 157085730, 109254766, 208403048, 237620966, 111341228, 210568560, 177255039,
              76642651, 41084242, 201062854, 130295133, 152865265, 175609590, 62045777, 118939950,
              168270865, 71471012, 235204060, 131798756, 162373432, 74680748, 112472991, 145384235}))
  stage_4_butterfly_6 (
    .x_in(stage_3_per_out[12]),
    .y_in(stage_3_per_out[13]),
    .x_out(stage_4_per_in[12]),
    .y_out(stage_4_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 197787791, 215696667, 172642311, 153962078, 11695616, 233560477, 189907315,
              181852808, 147699054, 146694818, 202366126, 218546733, 78852289, 227611463, 71460019,
              17079898, 193045667, 25574347, 66112528, 263678998, 115957373, 27685019, 47317233,
              179817683, 109553202, 6323336, 165226744, 200054106, 191662816, 170752771, 140204941,
              141548072, 169276669, 70982951, 119224607, 124918999, 82771912, 39593842, 239095400,
              102065274, 157085730, 109254766, 208403048, 237620966, 111341228, 210568560, 177255039,
              76642651, 41084242, 201062854, 130295133, 152865265, 175609590, 62045777, 118939950,
              168270865, 71471012, 235204060, 131798756, 162373432, 74680748, 112472991, 145384235}))
  stage_4_butterfly_7 (
    .x_in(stage_3_per_out[14]),
    .y_in(stage_3_per_out[15]),
    .x_out(stage_4_per_in[14]),
    .y_out(stage_4_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 197787791, 215696667, 172642311, 153962078, 11695616, 233560477, 189907315,
              181852808, 147699054, 146694818, 202366126, 218546733, 78852289, 227611463, 71460019,
              17079898, 193045667, 25574347, 66112528, 263678998, 115957373, 27685019, 47317233,
              179817683, 109553202, 6323336, 165226744, 200054106, 191662816, 170752771, 140204941,
              141548072, 169276669, 70982951, 119224607, 124918999, 82771912, 39593842, 239095400,
              102065274, 157085730, 109254766, 208403048, 237620966, 111341228, 210568560, 177255039,
              76642651, 41084242, 201062854, 130295133, 152865265, 175609590, 62045777, 118939950,
              168270865, 71471012, 235204060, 131798756, 162373432, 74680748, 112472991, 145384235}))
  stage_4_butterfly_8 (
    .x_in(stage_3_per_out[16]),
    .y_in(stage_3_per_out[17]),
    .x_out(stage_4_per_in[16]),
    .y_out(stage_4_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 197787791, 215696667, 172642311, 153962078, 11695616, 233560477, 189907315,
              181852808, 147699054, 146694818, 202366126, 218546733, 78852289, 227611463, 71460019,
              17079898, 193045667, 25574347, 66112528, 263678998, 115957373, 27685019, 47317233,
              179817683, 109553202, 6323336, 165226744, 200054106, 191662816, 170752771, 140204941,
              141548072, 169276669, 70982951, 119224607, 124918999, 82771912, 39593842, 239095400,
              102065274, 157085730, 109254766, 208403048, 237620966, 111341228, 210568560, 177255039,
              76642651, 41084242, 201062854, 130295133, 152865265, 175609590, 62045777, 118939950,
              168270865, 71471012, 235204060, 131798756, 162373432, 74680748, 112472991, 145384235}))
  stage_4_butterfly_9 (
    .x_in(stage_3_per_out[18]),
    .y_in(stage_3_per_out[19]),
    .x_out(stage_4_per_in[18]),
    .y_out(stage_4_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 197787791, 215696667, 172642311, 153962078, 11695616, 233560477, 189907315,
              181852808, 147699054, 146694818, 202366126, 218546733, 78852289, 227611463, 71460019,
              17079898, 193045667, 25574347, 66112528, 263678998, 115957373, 27685019, 47317233,
              179817683, 109553202, 6323336, 165226744, 200054106, 191662816, 170752771, 140204941,
              141548072, 169276669, 70982951, 119224607, 124918999, 82771912, 39593842, 239095400,
              102065274, 157085730, 109254766, 208403048, 237620966, 111341228, 210568560, 177255039,
              76642651, 41084242, 201062854, 130295133, 152865265, 175609590, 62045777, 118939950,
              168270865, 71471012, 235204060, 131798756, 162373432, 74680748, 112472991, 145384235}))
  stage_4_butterfly_10 (
    .x_in(stage_3_per_out[20]),
    .y_in(stage_3_per_out[21]),
    .x_out(stage_4_per_in[20]),
    .y_out(stage_4_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 197787791, 215696667, 172642311, 153962078, 11695616, 233560477, 189907315,
              181852808, 147699054, 146694818, 202366126, 218546733, 78852289, 227611463, 71460019,
              17079898, 193045667, 25574347, 66112528, 263678998, 115957373, 27685019, 47317233,
              179817683, 109553202, 6323336, 165226744, 200054106, 191662816, 170752771, 140204941,
              141548072, 169276669, 70982951, 119224607, 124918999, 82771912, 39593842, 239095400,
              102065274, 157085730, 109254766, 208403048, 237620966, 111341228, 210568560, 177255039,
              76642651, 41084242, 201062854, 130295133, 152865265, 175609590, 62045777, 118939950,
              168270865, 71471012, 235204060, 131798756, 162373432, 74680748, 112472991, 145384235}))
  stage_4_butterfly_11 (
    .x_in(stage_3_per_out[22]),
    .y_in(stage_3_per_out[23]),
    .x_out(stage_4_per_in[22]),
    .y_out(stage_4_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 197787791, 215696667, 172642311, 153962078, 11695616, 233560477, 189907315,
              181852808, 147699054, 146694818, 202366126, 218546733, 78852289, 227611463, 71460019,
              17079898, 193045667, 25574347, 66112528, 263678998, 115957373, 27685019, 47317233,
              179817683, 109553202, 6323336, 165226744, 200054106, 191662816, 170752771, 140204941,
              141548072, 169276669, 70982951, 119224607, 124918999, 82771912, 39593842, 239095400,
              102065274, 157085730, 109254766, 208403048, 237620966, 111341228, 210568560, 177255039,
              76642651, 41084242, 201062854, 130295133, 152865265, 175609590, 62045777, 118939950,
              168270865, 71471012, 235204060, 131798756, 162373432, 74680748, 112472991, 145384235}))
  stage_4_butterfly_12 (
    .x_in(stage_3_per_out[24]),
    .y_in(stage_3_per_out[25]),
    .x_out(stage_4_per_in[24]),
    .y_out(stage_4_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 197787791, 215696667, 172642311, 153962078, 11695616, 233560477, 189907315,
              181852808, 147699054, 146694818, 202366126, 218546733, 78852289, 227611463, 71460019,
              17079898, 193045667, 25574347, 66112528, 263678998, 115957373, 27685019, 47317233,
              179817683, 109553202, 6323336, 165226744, 200054106, 191662816, 170752771, 140204941,
              141548072, 169276669, 70982951, 119224607, 124918999, 82771912, 39593842, 239095400,
              102065274, 157085730, 109254766, 208403048, 237620966, 111341228, 210568560, 177255039,
              76642651, 41084242, 201062854, 130295133, 152865265, 175609590, 62045777, 118939950,
              168270865, 71471012, 235204060, 131798756, 162373432, 74680748, 112472991, 145384235}))
  stage_4_butterfly_13 (
    .x_in(stage_3_per_out[26]),
    .y_in(stage_3_per_out[27]),
    .x_out(stage_4_per_in[26]),
    .y_out(stage_4_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 197787791, 215696667, 172642311, 153962078, 11695616, 233560477, 189907315,
              181852808, 147699054, 146694818, 202366126, 218546733, 78852289, 227611463, 71460019,
              17079898, 193045667, 25574347, 66112528, 263678998, 115957373, 27685019, 47317233,
              179817683, 109553202, 6323336, 165226744, 200054106, 191662816, 170752771, 140204941,
              141548072, 169276669, 70982951, 119224607, 124918999, 82771912, 39593842, 239095400,
              102065274, 157085730, 109254766, 208403048, 237620966, 111341228, 210568560, 177255039,
              76642651, 41084242, 201062854, 130295133, 152865265, 175609590, 62045777, 118939950,
              168270865, 71471012, 235204060, 131798756, 162373432, 74680748, 112472991, 145384235}))
  stage_4_butterfly_14 (
    .x_in(stage_3_per_out[28]),
    .y_in(stage_3_per_out[29]),
    .x_out(stage_4_per_in[28]),
    .y_out(stage_4_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({92577793, 197787791, 215696667, 172642311, 153962078, 11695616, 233560477, 189907315,
              181852808, 147699054, 146694818, 202366126, 218546733, 78852289, 227611463, 71460019,
              17079898, 193045667, 25574347, 66112528, 263678998, 115957373, 27685019, 47317233,
              179817683, 109553202, 6323336, 165226744, 200054106, 191662816, 170752771, 140204941,
              141548072, 169276669, 70982951, 119224607, 124918999, 82771912, 39593842, 239095400,
              102065274, 157085730, 109254766, 208403048, 237620966, 111341228, 210568560, 177255039,
              76642651, 41084242, 201062854, 130295133, 152865265, 175609590, 62045777, 118939950,
              168270865, 71471012, 235204060, 131798756, 162373432, 74680748, 112472991, 145384235}))
  stage_4_butterfly_15 (
    .x_in(stage_3_per_out[30]),
    .y_in(stage_3_per_out[31]),
    .x_out(stage_4_per_in[30]),
    .y_out(stage_4_per_in[31]),
    .clk(clk),
    .rst(rst)
  );




  // TODO(Yang): stage 4 -> stage 5 permutation
  // FIXME: ignore butterfly units for now.
  stage_4_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_4_5_per (
    .inData_0(stage_4_per_in[0]),
    .inData_1(stage_4_per_in[1]),
    .inData_2(stage_4_per_in[2]),
    .inData_3(stage_4_per_in[3]),
    .inData_4(stage_4_per_in[4]),
    .inData_5(stage_4_per_in[5]),
    .inData_6(stage_4_per_in[6]),
    .inData_7(stage_4_per_in[7]),
    .inData_8(stage_4_per_in[8]),
    .inData_9(stage_4_per_in[9]),
    .inData_10(stage_4_per_in[10]),
    .inData_11(stage_4_per_in[11]),
    .inData_12(stage_4_per_in[12]),
    .inData_13(stage_4_per_in[13]),
    .inData_14(stage_4_per_in[14]),
    .inData_15(stage_4_per_in[15]),
    .inData_16(stage_4_per_in[16]),
    .inData_17(stage_4_per_in[17]),
    .inData_18(stage_4_per_in[18]),
    .inData_19(stage_4_per_in[19]),
    .inData_20(stage_4_per_in[20]),
    .inData_21(stage_4_per_in[21]),
    .inData_22(stage_4_per_in[22]),
    .inData_23(stage_4_per_in[23]),
    .inData_24(stage_4_per_in[24]),
    .inData_25(stage_4_per_in[25]),
    .inData_26(stage_4_per_in[26]),
    .inData_27(stage_4_per_in[27]),
    .inData_28(stage_4_per_in[28]),
    .inData_29(stage_4_per_in[29]),
    .inData_30(stage_4_per_in[30]),
    .inData_31(stage_4_per_in[31]),
    .outData_0(stage_4_per_out[0]),
    .outData_1(stage_4_per_out[1]),
    .outData_2(stage_4_per_out[2]),
    .outData_3(stage_4_per_out[3]),
    .outData_4(stage_4_per_out[4]),
    .outData_5(stage_4_per_out[5]),
    .outData_6(stage_4_per_out[6]),
    .outData_7(stage_4_per_out[7]),
    .outData_8(stage_4_per_out[8]),
    .outData_9(stage_4_per_out[9]),
    .outData_10(stage_4_per_out[10]),
    .outData_11(stage_4_per_out[11]),
    .outData_12(stage_4_per_out[12]),
    .outData_13(stage_4_per_out[13]),
    .outData_14(stage_4_per_out[14]),
    .outData_15(stage_4_per_out[15]),
    .outData_16(stage_4_per_out[16]),
    .outData_17(stage_4_per_out[17]),
    .outData_18(stage_4_per_out[18]),
    .outData_19(stage_4_per_out[19]),
    .outData_20(stage_4_per_out[20]),
    .outData_21(stage_4_per_out[21]),
    .outData_22(stage_4_per_out[22]),
    .outData_23(stage_4_per_out[23]),
    .outData_24(stage_4_per_out[24]),
    .outData_25(stage_4_per_out[25]),
    .outData_26(stage_4_per_out[26]),
    .outData_27(stage_4_per_out[27]),
    .outData_28(stage_4_per_out[28]),
    .outData_29(stage_4_per_out[29]),
    .outData_30(stage_4_per_out[30]),
    .outData_31(stage_4_per_out[31]),
    .in_start(in_start[4]),
    .out_start(out_start[4]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 5 32 butterfly units
  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 183300662, 108349160, 108349160, 178374402, 178374402, 220656190, 220656190,
              174234737, 174234737, 36955649, 36955649, 216372172, 216372172, 221840088, 221840088,
              249274747, 249274747, 206308099, 206308099, 35289455, 35289455, 76573097, 76573097,
              11699091, 11699091, 143639106, 143639106, 234642902, 234642902, 39264098, 39264098,
              57538295, 57538295, 84893967, 84893967, 265190919, 265190919, 165596304, 165596304,
              102579498, 102579498, 119480423, 119480423, 139368110, 139368110, 72061017, 72061017,
              92744225, 92744225, 5258704, 5258704, 83571649, 83571649, 220492738, 220492738,
              18533839, 18533839, 99790517, 99790517, 196317032, 196317032, 73825164, 73825164}))
  stage_5_butterfly_0 (
    .x_in(stage_4_per_out[0]),
    .y_in(stage_4_per_out[1]),
    .x_out(stage_5_per_in[0]),
    .y_out(stage_5_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 183300662, 108349160, 108349160, 178374402, 178374402, 220656190, 220656190,
              174234737, 174234737, 36955649, 36955649, 216372172, 216372172, 221840088, 221840088,
              249274747, 249274747, 206308099, 206308099, 35289455, 35289455, 76573097, 76573097,
              11699091, 11699091, 143639106, 143639106, 234642902, 234642902, 39264098, 39264098,
              57538295, 57538295, 84893967, 84893967, 265190919, 265190919, 165596304, 165596304,
              102579498, 102579498, 119480423, 119480423, 139368110, 139368110, 72061017, 72061017,
              92744225, 92744225, 5258704, 5258704, 83571649, 83571649, 220492738, 220492738,
              18533839, 18533839, 99790517, 99790517, 196317032, 196317032, 73825164, 73825164}))
  stage_5_butterfly_1 (
    .x_in(stage_4_per_out[2]),
    .y_in(stage_4_per_out[3]),
    .x_out(stage_5_per_in[2]),
    .y_out(stage_5_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 183300662, 108349160, 108349160, 178374402, 178374402, 220656190, 220656190,
              174234737, 174234737, 36955649, 36955649, 216372172, 216372172, 221840088, 221840088,
              249274747, 249274747, 206308099, 206308099, 35289455, 35289455, 76573097, 76573097,
              11699091, 11699091, 143639106, 143639106, 234642902, 234642902, 39264098, 39264098,
              57538295, 57538295, 84893967, 84893967, 265190919, 265190919, 165596304, 165596304,
              102579498, 102579498, 119480423, 119480423, 139368110, 139368110, 72061017, 72061017,
              92744225, 92744225, 5258704, 5258704, 83571649, 83571649, 220492738, 220492738,
              18533839, 18533839, 99790517, 99790517, 196317032, 196317032, 73825164, 73825164}))
  stage_5_butterfly_2 (
    .x_in(stage_4_per_out[4]),
    .y_in(stage_4_per_out[5]),
    .x_out(stage_5_per_in[4]),
    .y_out(stage_5_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 183300662, 108349160, 108349160, 178374402, 178374402, 220656190, 220656190,
              174234737, 174234737, 36955649, 36955649, 216372172, 216372172, 221840088, 221840088,
              249274747, 249274747, 206308099, 206308099, 35289455, 35289455, 76573097, 76573097,
              11699091, 11699091, 143639106, 143639106, 234642902, 234642902, 39264098, 39264098,
              57538295, 57538295, 84893967, 84893967, 265190919, 265190919, 165596304, 165596304,
              102579498, 102579498, 119480423, 119480423, 139368110, 139368110, 72061017, 72061017,
              92744225, 92744225, 5258704, 5258704, 83571649, 83571649, 220492738, 220492738,
              18533839, 18533839, 99790517, 99790517, 196317032, 196317032, 73825164, 73825164}))
  stage_5_butterfly_3 (
    .x_in(stage_4_per_out[6]),
    .y_in(stage_4_per_out[7]),
    .x_out(stage_5_per_in[6]),
    .y_out(stage_5_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 183300662, 108349160, 108349160, 178374402, 178374402, 220656190, 220656190,
              174234737, 174234737, 36955649, 36955649, 216372172, 216372172, 221840088, 221840088,
              249274747, 249274747, 206308099, 206308099, 35289455, 35289455, 76573097, 76573097,
              11699091, 11699091, 143639106, 143639106, 234642902, 234642902, 39264098, 39264098,
              57538295, 57538295, 84893967, 84893967, 265190919, 265190919, 165596304, 165596304,
              102579498, 102579498, 119480423, 119480423, 139368110, 139368110, 72061017, 72061017,
              92744225, 92744225, 5258704, 5258704, 83571649, 83571649, 220492738, 220492738,
              18533839, 18533839, 99790517, 99790517, 196317032, 196317032, 73825164, 73825164}))
  stage_5_butterfly_4 (
    .x_in(stage_4_per_out[8]),
    .y_in(stage_4_per_out[9]),
    .x_out(stage_5_per_in[8]),
    .y_out(stage_5_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 183300662, 108349160, 108349160, 178374402, 178374402, 220656190, 220656190,
              174234737, 174234737, 36955649, 36955649, 216372172, 216372172, 221840088, 221840088,
              249274747, 249274747, 206308099, 206308099, 35289455, 35289455, 76573097, 76573097,
              11699091, 11699091, 143639106, 143639106, 234642902, 234642902, 39264098, 39264098,
              57538295, 57538295, 84893967, 84893967, 265190919, 265190919, 165596304, 165596304,
              102579498, 102579498, 119480423, 119480423, 139368110, 139368110, 72061017, 72061017,
              92744225, 92744225, 5258704, 5258704, 83571649, 83571649, 220492738, 220492738,
              18533839, 18533839, 99790517, 99790517, 196317032, 196317032, 73825164, 73825164}))
  stage_5_butterfly_5 (
    .x_in(stage_4_per_out[10]),
    .y_in(stage_4_per_out[11]),
    .x_out(stage_5_per_in[10]),
    .y_out(stage_5_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 183300662, 108349160, 108349160, 178374402, 178374402, 220656190, 220656190,
              174234737, 174234737, 36955649, 36955649, 216372172, 216372172, 221840088, 221840088,
              249274747, 249274747, 206308099, 206308099, 35289455, 35289455, 76573097, 76573097,
              11699091, 11699091, 143639106, 143639106, 234642902, 234642902, 39264098, 39264098,
              57538295, 57538295, 84893967, 84893967, 265190919, 265190919, 165596304, 165596304,
              102579498, 102579498, 119480423, 119480423, 139368110, 139368110, 72061017, 72061017,
              92744225, 92744225, 5258704, 5258704, 83571649, 83571649, 220492738, 220492738,
              18533839, 18533839, 99790517, 99790517, 196317032, 196317032, 73825164, 73825164}))
  stage_5_butterfly_6 (
    .x_in(stage_4_per_out[12]),
    .y_in(stage_4_per_out[13]),
    .x_out(stage_5_per_in[12]),
    .y_out(stage_5_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 183300662, 108349160, 108349160, 178374402, 178374402, 220656190, 220656190,
              174234737, 174234737, 36955649, 36955649, 216372172, 216372172, 221840088, 221840088,
              249274747, 249274747, 206308099, 206308099, 35289455, 35289455, 76573097, 76573097,
              11699091, 11699091, 143639106, 143639106, 234642902, 234642902, 39264098, 39264098,
              57538295, 57538295, 84893967, 84893967, 265190919, 265190919, 165596304, 165596304,
              102579498, 102579498, 119480423, 119480423, 139368110, 139368110, 72061017, 72061017,
              92744225, 92744225, 5258704, 5258704, 83571649, 83571649, 220492738, 220492738,
              18533839, 18533839, 99790517, 99790517, 196317032, 196317032, 73825164, 73825164}))
  stage_5_butterfly_7 (
    .x_in(stage_4_per_out[14]),
    .y_in(stage_4_per_out[15]),
    .x_out(stage_5_per_in[14]),
    .y_out(stage_5_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 183300662, 108349160, 108349160, 178374402, 178374402, 220656190, 220656190,
              174234737, 174234737, 36955649, 36955649, 216372172, 216372172, 221840088, 221840088,
              249274747, 249274747, 206308099, 206308099, 35289455, 35289455, 76573097, 76573097,
              11699091, 11699091, 143639106, 143639106, 234642902, 234642902, 39264098, 39264098,
              57538295, 57538295, 84893967, 84893967, 265190919, 265190919, 165596304, 165596304,
              102579498, 102579498, 119480423, 119480423, 139368110, 139368110, 72061017, 72061017,
              92744225, 92744225, 5258704, 5258704, 83571649, 83571649, 220492738, 220492738,
              18533839, 18533839, 99790517, 99790517, 196317032, 196317032, 73825164, 73825164}))
  stage_5_butterfly_8 (
    .x_in(stage_4_per_out[16]),
    .y_in(stage_4_per_out[17]),
    .x_out(stage_5_per_in[16]),
    .y_out(stage_5_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 183300662, 108349160, 108349160, 178374402, 178374402, 220656190, 220656190,
              174234737, 174234737, 36955649, 36955649, 216372172, 216372172, 221840088, 221840088,
              249274747, 249274747, 206308099, 206308099, 35289455, 35289455, 76573097, 76573097,
              11699091, 11699091, 143639106, 143639106, 234642902, 234642902, 39264098, 39264098,
              57538295, 57538295, 84893967, 84893967, 265190919, 265190919, 165596304, 165596304,
              102579498, 102579498, 119480423, 119480423, 139368110, 139368110, 72061017, 72061017,
              92744225, 92744225, 5258704, 5258704, 83571649, 83571649, 220492738, 220492738,
              18533839, 18533839, 99790517, 99790517, 196317032, 196317032, 73825164, 73825164}))
  stage_5_butterfly_9 (
    .x_in(stage_4_per_out[18]),
    .y_in(stage_4_per_out[19]),
    .x_out(stage_5_per_in[18]),
    .y_out(stage_5_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 183300662, 108349160, 108349160, 178374402, 178374402, 220656190, 220656190,
              174234737, 174234737, 36955649, 36955649, 216372172, 216372172, 221840088, 221840088,
              249274747, 249274747, 206308099, 206308099, 35289455, 35289455, 76573097, 76573097,
              11699091, 11699091, 143639106, 143639106, 234642902, 234642902, 39264098, 39264098,
              57538295, 57538295, 84893967, 84893967, 265190919, 265190919, 165596304, 165596304,
              102579498, 102579498, 119480423, 119480423, 139368110, 139368110, 72061017, 72061017,
              92744225, 92744225, 5258704, 5258704, 83571649, 83571649, 220492738, 220492738,
              18533839, 18533839, 99790517, 99790517, 196317032, 196317032, 73825164, 73825164}))
  stage_5_butterfly_10 (
    .x_in(stage_4_per_out[20]),
    .y_in(stage_4_per_out[21]),
    .x_out(stage_5_per_in[20]),
    .y_out(stage_5_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 183300662, 108349160, 108349160, 178374402, 178374402, 220656190, 220656190,
              174234737, 174234737, 36955649, 36955649, 216372172, 216372172, 221840088, 221840088,
              249274747, 249274747, 206308099, 206308099, 35289455, 35289455, 76573097, 76573097,
              11699091, 11699091, 143639106, 143639106, 234642902, 234642902, 39264098, 39264098,
              57538295, 57538295, 84893967, 84893967, 265190919, 265190919, 165596304, 165596304,
              102579498, 102579498, 119480423, 119480423, 139368110, 139368110, 72061017, 72061017,
              92744225, 92744225, 5258704, 5258704, 83571649, 83571649, 220492738, 220492738,
              18533839, 18533839, 99790517, 99790517, 196317032, 196317032, 73825164, 73825164}))
  stage_5_butterfly_11 (
    .x_in(stage_4_per_out[22]),
    .y_in(stage_4_per_out[23]),
    .x_out(stage_5_per_in[22]),
    .y_out(stage_5_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 183300662, 108349160, 108349160, 178374402, 178374402, 220656190, 220656190,
              174234737, 174234737, 36955649, 36955649, 216372172, 216372172, 221840088, 221840088,
              249274747, 249274747, 206308099, 206308099, 35289455, 35289455, 76573097, 76573097,
              11699091, 11699091, 143639106, 143639106, 234642902, 234642902, 39264098, 39264098,
              57538295, 57538295, 84893967, 84893967, 265190919, 265190919, 165596304, 165596304,
              102579498, 102579498, 119480423, 119480423, 139368110, 139368110, 72061017, 72061017,
              92744225, 92744225, 5258704, 5258704, 83571649, 83571649, 220492738, 220492738,
              18533839, 18533839, 99790517, 99790517, 196317032, 196317032, 73825164, 73825164}))
  stage_5_butterfly_12 (
    .x_in(stage_4_per_out[24]),
    .y_in(stage_4_per_out[25]),
    .x_out(stage_5_per_in[24]),
    .y_out(stage_5_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 183300662, 108349160, 108349160, 178374402, 178374402, 220656190, 220656190,
              174234737, 174234737, 36955649, 36955649, 216372172, 216372172, 221840088, 221840088,
              249274747, 249274747, 206308099, 206308099, 35289455, 35289455, 76573097, 76573097,
              11699091, 11699091, 143639106, 143639106, 234642902, 234642902, 39264098, 39264098,
              57538295, 57538295, 84893967, 84893967, 265190919, 265190919, 165596304, 165596304,
              102579498, 102579498, 119480423, 119480423, 139368110, 139368110, 72061017, 72061017,
              92744225, 92744225, 5258704, 5258704, 83571649, 83571649, 220492738, 220492738,
              18533839, 18533839, 99790517, 99790517, 196317032, 196317032, 73825164, 73825164}))
  stage_5_butterfly_13 (
    .x_in(stage_4_per_out[26]),
    .y_in(stage_4_per_out[27]),
    .x_out(stage_5_per_in[26]),
    .y_out(stage_5_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 183300662, 108349160, 108349160, 178374402, 178374402, 220656190, 220656190,
              174234737, 174234737, 36955649, 36955649, 216372172, 216372172, 221840088, 221840088,
              249274747, 249274747, 206308099, 206308099, 35289455, 35289455, 76573097, 76573097,
              11699091, 11699091, 143639106, 143639106, 234642902, 234642902, 39264098, 39264098,
              57538295, 57538295, 84893967, 84893967, 265190919, 265190919, 165596304, 165596304,
              102579498, 102579498, 119480423, 119480423, 139368110, 139368110, 72061017, 72061017,
              92744225, 92744225, 5258704, 5258704, 83571649, 83571649, 220492738, 220492738,
              18533839, 18533839, 99790517, 99790517, 196317032, 196317032, 73825164, 73825164}))
  stage_5_butterfly_14 (
    .x_in(stage_4_per_out[28]),
    .y_in(stage_4_per_out[29]),
    .x_out(stage_5_per_in[28]),
    .y_out(stage_5_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({183300662, 183300662, 108349160, 108349160, 178374402, 178374402, 220656190, 220656190,
              174234737, 174234737, 36955649, 36955649, 216372172, 216372172, 221840088, 221840088,
              249274747, 249274747, 206308099, 206308099, 35289455, 35289455, 76573097, 76573097,
              11699091, 11699091, 143639106, 143639106, 234642902, 234642902, 39264098, 39264098,
              57538295, 57538295, 84893967, 84893967, 265190919, 265190919, 165596304, 165596304,
              102579498, 102579498, 119480423, 119480423, 139368110, 139368110, 72061017, 72061017,
              92744225, 92744225, 5258704, 5258704, 83571649, 83571649, 220492738, 220492738,
              18533839, 18533839, 99790517, 99790517, 196317032, 196317032, 73825164, 73825164}))
  stage_5_butterfly_15 (
    .x_in(stage_4_per_out[30]),
    .y_in(stage_4_per_out[31]),
    .x_out(stage_5_per_in[30]),
    .y_out(stage_5_per_in[31]),
    .clk(clk),
    .rst(rst)
  );





  // TODO(Yang): stage 5 -> stage 6 permutation
  // FIXME: ignore butterfly units for now.
  stage_5_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_5_6_per (
    .inData_0(stage_5_per_in[0]),
    .inData_1(stage_5_per_in[1]),
    .inData_2(stage_5_per_in[2]),
    .inData_3(stage_5_per_in[3]),
    .inData_4(stage_5_per_in[4]),
    .inData_5(stage_5_per_in[5]),
    .inData_6(stage_5_per_in[6]),
    .inData_7(stage_5_per_in[7]),
    .inData_8(stage_5_per_in[8]),
    .inData_9(stage_5_per_in[9]),
    .inData_10(stage_5_per_in[10]),
    .inData_11(stage_5_per_in[11]),
    .inData_12(stage_5_per_in[12]),
    .inData_13(stage_5_per_in[13]),
    .inData_14(stage_5_per_in[14]),
    .inData_15(stage_5_per_in[15]),
    .inData_16(stage_5_per_in[16]),
    .inData_17(stage_5_per_in[17]),
    .inData_18(stage_5_per_in[18]),
    .inData_19(stage_5_per_in[19]),
    .inData_20(stage_5_per_in[20]),
    .inData_21(stage_5_per_in[21]),
    .inData_22(stage_5_per_in[22]),
    .inData_23(stage_5_per_in[23]),
    .inData_24(stage_5_per_in[24]),
    .inData_25(stage_5_per_in[25]),
    .inData_26(stage_5_per_in[26]),
    .inData_27(stage_5_per_in[27]),
    .inData_28(stage_5_per_in[28]),
    .inData_29(stage_5_per_in[29]),
    .inData_30(stage_5_per_in[30]),
    .inData_31(stage_5_per_in[31]),
    .outData_0(stage_5_per_out[0]),
    .outData_1(stage_5_per_out[1]),
    .outData_2(stage_5_per_out[2]),
    .outData_3(stage_5_per_out[3]),
    .outData_4(stage_5_per_out[4]),
    .outData_5(stage_5_per_out[5]),
    .outData_6(stage_5_per_out[6]),
    .outData_7(stage_5_per_out[7]),
    .outData_8(stage_5_per_out[8]),
    .outData_9(stage_5_per_out[9]),
    .outData_10(stage_5_per_out[10]),
    .outData_11(stage_5_per_out[11]),
    .outData_12(stage_5_per_out[12]),
    .outData_13(stage_5_per_out[13]),
    .outData_14(stage_5_per_out[14]),
    .outData_15(stage_5_per_out[15]),
    .outData_16(stage_5_per_out[16]),
    .outData_17(stage_5_per_out[17]),
    .outData_18(stage_5_per_out[18]),
    .outData_19(stage_5_per_out[19]),
    .outData_20(stage_5_per_out[20]),
    .outData_21(stage_5_per_out[21]),
    .outData_22(stage_5_per_out[22]),
    .outData_23(stage_5_per_out[23]),
    .outData_24(stage_5_per_out[24]),
    .outData_25(stage_5_per_out[25]),
    .outData_26(stage_5_per_out[26]),
    .outData_27(stage_5_per_out[27]),
    .outData_28(stage_5_per_out[28]),
    .outData_29(stage_5_per_out[29]),
    .outData_30(stage_5_per_out[30]),
    .outData_31(stage_5_per_out[31]),
    .in_start(in_start[5]),
    .out_start(out_start[5]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 6 32 butterfly units
  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 73648196, 73648196, 163057267, 163057267, 163057267, 163057267,
              42982065, 42982065, 42982065, 42982065, 135333989, 135333989, 135333989, 135333989,
              46265048, 46265048, 46265048, 46265048, 242569099, 242569099, 242569099, 242569099,
              70516281, 70516281, 70516281, 70516281, 136955445, 136955445, 136955445, 136955445,
              33383981, 33383981, 33383981, 33383981, 47600907, 47600907, 47600907, 47600907,
              142393906, 142393906, 142393906, 142393906, 69075086, 69075086, 69075086, 69075086,
              210749829, 210749829, 210749829, 210749829, 133782759, 133782759, 133782759, 133782759,
              155624840, 155624840, 155624840, 155624840, 7802111, 7802111, 7802111, 7802111}))
  stage_6_butterfly_0 (
    .x_in(stage_5_per_out[0]),
    .y_in(stage_5_per_out[1]),
    .x_out(stage_6_per_in[0]),
    .y_out(stage_6_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 73648196, 73648196, 163057267, 163057267, 163057267, 163057267,
              42982065, 42982065, 42982065, 42982065, 135333989, 135333989, 135333989, 135333989,
              46265048, 46265048, 46265048, 46265048, 242569099, 242569099, 242569099, 242569099,
              70516281, 70516281, 70516281, 70516281, 136955445, 136955445, 136955445, 136955445,
              33383981, 33383981, 33383981, 33383981, 47600907, 47600907, 47600907, 47600907,
              142393906, 142393906, 142393906, 142393906, 69075086, 69075086, 69075086, 69075086,
              210749829, 210749829, 210749829, 210749829, 133782759, 133782759, 133782759, 133782759,
              155624840, 155624840, 155624840, 155624840, 7802111, 7802111, 7802111, 7802111}))
  stage_6_butterfly_1 (
    .x_in(stage_5_per_out[2]),
    .y_in(stage_5_per_out[3]),
    .x_out(stage_6_per_in[2]),
    .y_out(stage_6_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 73648196, 73648196, 163057267, 163057267, 163057267, 163057267,
              42982065, 42982065, 42982065, 42982065, 135333989, 135333989, 135333989, 135333989,
              46265048, 46265048, 46265048, 46265048, 242569099, 242569099, 242569099, 242569099,
              70516281, 70516281, 70516281, 70516281, 136955445, 136955445, 136955445, 136955445,
              33383981, 33383981, 33383981, 33383981, 47600907, 47600907, 47600907, 47600907,
              142393906, 142393906, 142393906, 142393906, 69075086, 69075086, 69075086, 69075086,
              210749829, 210749829, 210749829, 210749829, 133782759, 133782759, 133782759, 133782759,
              155624840, 155624840, 155624840, 155624840, 7802111, 7802111, 7802111, 7802111}))
  stage_6_butterfly_2 (
    .x_in(stage_5_per_out[4]),
    .y_in(stage_5_per_out[5]),
    .x_out(stage_6_per_in[4]),
    .y_out(stage_6_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 73648196, 73648196, 163057267, 163057267, 163057267, 163057267,
              42982065, 42982065, 42982065, 42982065, 135333989, 135333989, 135333989, 135333989,
              46265048, 46265048, 46265048, 46265048, 242569099, 242569099, 242569099, 242569099,
              70516281, 70516281, 70516281, 70516281, 136955445, 136955445, 136955445, 136955445,
              33383981, 33383981, 33383981, 33383981, 47600907, 47600907, 47600907, 47600907,
              142393906, 142393906, 142393906, 142393906, 69075086, 69075086, 69075086, 69075086,
              210749829, 210749829, 210749829, 210749829, 133782759, 133782759, 133782759, 133782759,
              155624840, 155624840, 155624840, 155624840, 7802111, 7802111, 7802111, 7802111}))
  stage_6_butterfly_3 (
    .x_in(stage_5_per_out[6]),
    .y_in(stage_5_per_out[7]),
    .x_out(stage_6_per_in[6]),
    .y_out(stage_6_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 73648196, 73648196, 163057267, 163057267, 163057267, 163057267,
              42982065, 42982065, 42982065, 42982065, 135333989, 135333989, 135333989, 135333989,
              46265048, 46265048, 46265048, 46265048, 242569099, 242569099, 242569099, 242569099,
              70516281, 70516281, 70516281, 70516281, 136955445, 136955445, 136955445, 136955445,
              33383981, 33383981, 33383981, 33383981, 47600907, 47600907, 47600907, 47600907,
              142393906, 142393906, 142393906, 142393906, 69075086, 69075086, 69075086, 69075086,
              210749829, 210749829, 210749829, 210749829, 133782759, 133782759, 133782759, 133782759,
              155624840, 155624840, 155624840, 155624840, 7802111, 7802111, 7802111, 7802111}))
  stage_6_butterfly_4 (
    .x_in(stage_5_per_out[8]),
    .y_in(stage_5_per_out[9]),
    .x_out(stage_6_per_in[8]),
    .y_out(stage_6_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 73648196, 73648196, 163057267, 163057267, 163057267, 163057267,
              42982065, 42982065, 42982065, 42982065, 135333989, 135333989, 135333989, 135333989,
              46265048, 46265048, 46265048, 46265048, 242569099, 242569099, 242569099, 242569099,
              70516281, 70516281, 70516281, 70516281, 136955445, 136955445, 136955445, 136955445,
              33383981, 33383981, 33383981, 33383981, 47600907, 47600907, 47600907, 47600907,
              142393906, 142393906, 142393906, 142393906, 69075086, 69075086, 69075086, 69075086,
              210749829, 210749829, 210749829, 210749829, 133782759, 133782759, 133782759, 133782759,
              155624840, 155624840, 155624840, 155624840, 7802111, 7802111, 7802111, 7802111}))
  stage_6_butterfly_5 (
    .x_in(stage_5_per_out[10]),
    .y_in(stage_5_per_out[11]),
    .x_out(stage_6_per_in[10]),
    .y_out(stage_6_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 73648196, 73648196, 163057267, 163057267, 163057267, 163057267,
              42982065, 42982065, 42982065, 42982065, 135333989, 135333989, 135333989, 135333989,
              46265048, 46265048, 46265048, 46265048, 242569099, 242569099, 242569099, 242569099,
              70516281, 70516281, 70516281, 70516281, 136955445, 136955445, 136955445, 136955445,
              33383981, 33383981, 33383981, 33383981, 47600907, 47600907, 47600907, 47600907,
              142393906, 142393906, 142393906, 142393906, 69075086, 69075086, 69075086, 69075086,
              210749829, 210749829, 210749829, 210749829, 133782759, 133782759, 133782759, 133782759,
              155624840, 155624840, 155624840, 155624840, 7802111, 7802111, 7802111, 7802111}))
  stage_6_butterfly_6 (
    .x_in(stage_5_per_out[12]),
    .y_in(stage_5_per_out[13]),
    .x_out(stage_6_per_in[12]),
    .y_out(stage_6_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 73648196, 73648196, 163057267, 163057267, 163057267, 163057267,
              42982065, 42982065, 42982065, 42982065, 135333989, 135333989, 135333989, 135333989,
              46265048, 46265048, 46265048, 46265048, 242569099, 242569099, 242569099, 242569099,
              70516281, 70516281, 70516281, 70516281, 136955445, 136955445, 136955445, 136955445,
              33383981, 33383981, 33383981, 33383981, 47600907, 47600907, 47600907, 47600907,
              142393906, 142393906, 142393906, 142393906, 69075086, 69075086, 69075086, 69075086,
              210749829, 210749829, 210749829, 210749829, 133782759, 133782759, 133782759, 133782759,
              155624840, 155624840, 155624840, 155624840, 7802111, 7802111, 7802111, 7802111}))
  stage_6_butterfly_7 (
    .x_in(stage_5_per_out[14]),
    .y_in(stage_5_per_out[15]),
    .x_out(stage_6_per_in[14]),
    .y_out(stage_6_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 73648196, 73648196, 163057267, 163057267, 163057267, 163057267,
              42982065, 42982065, 42982065, 42982065, 135333989, 135333989, 135333989, 135333989,
              46265048, 46265048, 46265048, 46265048, 242569099, 242569099, 242569099, 242569099,
              70516281, 70516281, 70516281, 70516281, 136955445, 136955445, 136955445, 136955445,
              33383981, 33383981, 33383981, 33383981, 47600907, 47600907, 47600907, 47600907,
              142393906, 142393906, 142393906, 142393906, 69075086, 69075086, 69075086, 69075086,
              210749829, 210749829, 210749829, 210749829, 133782759, 133782759, 133782759, 133782759,
              155624840, 155624840, 155624840, 155624840, 7802111, 7802111, 7802111, 7802111}))
  stage_6_butterfly_8 (
    .x_in(stage_5_per_out[16]),
    .y_in(stage_5_per_out[17]),
    .x_out(stage_6_per_in[16]),
    .y_out(stage_6_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 73648196, 73648196, 163057267, 163057267, 163057267, 163057267,
              42982065, 42982065, 42982065, 42982065, 135333989, 135333989, 135333989, 135333989,
              46265048, 46265048, 46265048, 46265048, 242569099, 242569099, 242569099, 242569099,
              70516281, 70516281, 70516281, 70516281, 136955445, 136955445, 136955445, 136955445,
              33383981, 33383981, 33383981, 33383981, 47600907, 47600907, 47600907, 47600907,
              142393906, 142393906, 142393906, 142393906, 69075086, 69075086, 69075086, 69075086,
              210749829, 210749829, 210749829, 210749829, 133782759, 133782759, 133782759, 133782759,
              155624840, 155624840, 155624840, 155624840, 7802111, 7802111, 7802111, 7802111}))
  stage_6_butterfly_9 (
    .x_in(stage_5_per_out[18]),
    .y_in(stage_5_per_out[19]),
    .x_out(stage_6_per_in[18]),
    .y_out(stage_6_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 73648196, 73648196, 163057267, 163057267, 163057267, 163057267,
              42982065, 42982065, 42982065, 42982065, 135333989, 135333989, 135333989, 135333989,
              46265048, 46265048, 46265048, 46265048, 242569099, 242569099, 242569099, 242569099,
              70516281, 70516281, 70516281, 70516281, 136955445, 136955445, 136955445, 136955445,
              33383981, 33383981, 33383981, 33383981, 47600907, 47600907, 47600907, 47600907,
              142393906, 142393906, 142393906, 142393906, 69075086, 69075086, 69075086, 69075086,
              210749829, 210749829, 210749829, 210749829, 133782759, 133782759, 133782759, 133782759,
              155624840, 155624840, 155624840, 155624840, 7802111, 7802111, 7802111, 7802111}))
  stage_6_butterfly_10 (
    .x_in(stage_5_per_out[20]),
    .y_in(stage_5_per_out[21]),
    .x_out(stage_6_per_in[20]),
    .y_out(stage_6_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 73648196, 73648196, 163057267, 163057267, 163057267, 163057267,
              42982065, 42982065, 42982065, 42982065, 135333989, 135333989, 135333989, 135333989,
              46265048, 46265048, 46265048, 46265048, 242569099, 242569099, 242569099, 242569099,
              70516281, 70516281, 70516281, 70516281, 136955445, 136955445, 136955445, 136955445,
              33383981, 33383981, 33383981, 33383981, 47600907, 47600907, 47600907, 47600907,
              142393906, 142393906, 142393906, 142393906, 69075086, 69075086, 69075086, 69075086,
              210749829, 210749829, 210749829, 210749829, 133782759, 133782759, 133782759, 133782759,
              155624840, 155624840, 155624840, 155624840, 7802111, 7802111, 7802111, 7802111}))
  stage_6_butterfly_11 (
    .x_in(stage_5_per_out[22]),
    .y_in(stage_5_per_out[23]),
    .x_out(stage_6_per_in[22]),
    .y_out(stage_6_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 73648196, 73648196, 163057267, 163057267, 163057267, 163057267,
              42982065, 42982065, 42982065, 42982065, 135333989, 135333989, 135333989, 135333989,
              46265048, 46265048, 46265048, 46265048, 242569099, 242569099, 242569099, 242569099,
              70516281, 70516281, 70516281, 70516281, 136955445, 136955445, 136955445, 136955445,
              33383981, 33383981, 33383981, 33383981, 47600907, 47600907, 47600907, 47600907,
              142393906, 142393906, 142393906, 142393906, 69075086, 69075086, 69075086, 69075086,
              210749829, 210749829, 210749829, 210749829, 133782759, 133782759, 133782759, 133782759,
              155624840, 155624840, 155624840, 155624840, 7802111, 7802111, 7802111, 7802111}))
  stage_6_butterfly_12 (
    .x_in(stage_5_per_out[24]),
    .y_in(stage_5_per_out[25]),
    .x_out(stage_6_per_in[24]),
    .y_out(stage_6_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 73648196, 73648196, 163057267, 163057267, 163057267, 163057267,
              42982065, 42982065, 42982065, 42982065, 135333989, 135333989, 135333989, 135333989,
              46265048, 46265048, 46265048, 46265048, 242569099, 242569099, 242569099, 242569099,
              70516281, 70516281, 70516281, 70516281, 136955445, 136955445, 136955445, 136955445,
              33383981, 33383981, 33383981, 33383981, 47600907, 47600907, 47600907, 47600907,
              142393906, 142393906, 142393906, 142393906, 69075086, 69075086, 69075086, 69075086,
              210749829, 210749829, 210749829, 210749829, 133782759, 133782759, 133782759, 133782759,
              155624840, 155624840, 155624840, 155624840, 7802111, 7802111, 7802111, 7802111}))
  stage_6_butterfly_13 (
    .x_in(stage_5_per_out[26]),
    .y_in(stage_5_per_out[27]),
    .x_out(stage_6_per_in[26]),
    .y_out(stage_6_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 73648196, 73648196, 163057267, 163057267, 163057267, 163057267,
              42982065, 42982065, 42982065, 42982065, 135333989, 135333989, 135333989, 135333989,
              46265048, 46265048, 46265048, 46265048, 242569099, 242569099, 242569099, 242569099,
              70516281, 70516281, 70516281, 70516281, 136955445, 136955445, 136955445, 136955445,
              33383981, 33383981, 33383981, 33383981, 47600907, 47600907, 47600907, 47600907,
              142393906, 142393906, 142393906, 142393906, 69075086, 69075086, 69075086, 69075086,
              210749829, 210749829, 210749829, 210749829, 133782759, 133782759, 133782759, 133782759,
              155624840, 155624840, 155624840, 155624840, 7802111, 7802111, 7802111, 7802111}))
  stage_6_butterfly_14 (
    .x_in(stage_5_per_out[28]),
    .y_in(stage_5_per_out[29]),
    .x_out(stage_6_per_in[28]),
    .y_out(stage_6_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({73648196, 73648196, 73648196, 73648196, 163057267, 163057267, 163057267, 163057267,
              42982065, 42982065, 42982065, 42982065, 135333989, 135333989, 135333989, 135333989,
              46265048, 46265048, 46265048, 46265048, 242569099, 242569099, 242569099, 242569099,
              70516281, 70516281, 70516281, 70516281, 136955445, 136955445, 136955445, 136955445,
              33383981, 33383981, 33383981, 33383981, 47600907, 47600907, 47600907, 47600907,
              142393906, 142393906, 142393906, 142393906, 69075086, 69075086, 69075086, 69075086,
              210749829, 210749829, 210749829, 210749829, 133782759, 133782759, 133782759, 133782759,
              155624840, 155624840, 155624840, 155624840, 7802111, 7802111, 7802111, 7802111}))
  stage_6_butterfly_15 (
    .x_in(stage_5_per_out[30]),
    .y_in(stage_5_per_out[31]),
    .x_out(stage_6_per_in[30]),
    .y_out(stage_6_per_in[31]),
    .clk(clk),
    .rst(rst)
  );




  // TODO(Yang): stage 6 -> stage 7 permutation
  // FIXME: ignore butterfly units for now.
  stage_6_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_6_7_per (
    .inData_0(stage_6_per_in[0]),
    .inData_1(stage_6_per_in[1]),
    .inData_2(stage_6_per_in[2]),
    .inData_3(stage_6_per_in[3]),
    .inData_4(stage_6_per_in[4]),
    .inData_5(stage_6_per_in[5]),
    .inData_6(stage_6_per_in[6]),
    .inData_7(stage_6_per_in[7]),
    .inData_8(stage_6_per_in[8]),
    .inData_9(stage_6_per_in[9]),
    .inData_10(stage_6_per_in[10]),
    .inData_11(stage_6_per_in[11]),
    .inData_12(stage_6_per_in[12]),
    .inData_13(stage_6_per_in[13]),
    .inData_14(stage_6_per_in[14]),
    .inData_15(stage_6_per_in[15]),
    .inData_16(stage_6_per_in[16]),
    .inData_17(stage_6_per_in[17]),
    .inData_18(stage_6_per_in[18]),
    .inData_19(stage_6_per_in[19]),
    .inData_20(stage_6_per_in[20]),
    .inData_21(stage_6_per_in[21]),
    .inData_22(stage_6_per_in[22]),
    .inData_23(stage_6_per_in[23]),
    .inData_24(stage_6_per_in[24]),
    .inData_25(stage_6_per_in[25]),
    .inData_26(stage_6_per_in[26]),
    .inData_27(stage_6_per_in[27]),
    .inData_28(stage_6_per_in[28]),
    .inData_29(stage_6_per_in[29]),
    .inData_30(stage_6_per_in[30]),
    .inData_31(stage_6_per_in[31]),
    .outData_0(stage_6_per_out[0]),
    .outData_1(stage_6_per_out[1]),
    .outData_2(stage_6_per_out[2]),
    .outData_3(stage_6_per_out[3]),
    .outData_4(stage_6_per_out[4]),
    .outData_5(stage_6_per_out[5]),
    .outData_6(stage_6_per_out[6]),
    .outData_7(stage_6_per_out[7]),
    .outData_8(stage_6_per_out[8]),
    .outData_9(stage_6_per_out[9]),
    .outData_10(stage_6_per_out[10]),
    .outData_11(stage_6_per_out[11]),
    .outData_12(stage_6_per_out[12]),
    .outData_13(stage_6_per_out[13]),
    .outData_14(stage_6_per_out[14]),
    .outData_15(stage_6_per_out[15]),
    .outData_16(stage_6_per_out[16]),
    .outData_17(stage_6_per_out[17]),
    .outData_18(stage_6_per_out[18]),
    .outData_19(stage_6_per_out[19]),
    .outData_20(stage_6_per_out[20]),
    .outData_21(stage_6_per_out[21]),
    .outData_22(stage_6_per_out[22]),
    .outData_23(stage_6_per_out[23]),
    .outData_24(stage_6_per_out[24]),
    .outData_25(stage_6_per_out[25]),
    .outData_26(stage_6_per_out[26]),
    .outData_27(stage_6_per_out[27]),
    .outData_28(stage_6_per_out[28]),
    .outData_29(stage_6_per_out[29]),
    .outData_30(stage_6_per_out[30]),
    .outData_31(stage_6_per_out[31]),
    .in_start(in_start[6]),
    .out_start(out_start[6]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 7 32 butterfly units
  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896,
              180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241,
              71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_0 (
    .x_in(stage_6_per_out[0]),
    .y_in(stage_6_per_out[1]),
    .x_out(stage_7_per_in[0]),
    .y_out(stage_7_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896,
              180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241,
              71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_1 (
    .x_in(stage_6_per_out[2]),
    .y_in(stage_6_per_out[3]),
    .x_out(stage_7_per_in[2]),
    .y_out(stage_7_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896,
              180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241,
              71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_2 (
    .x_in(stage_6_per_out[4]),
    .y_in(stage_6_per_out[5]),
    .x_out(stage_7_per_in[4]),
    .y_out(stage_7_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896,
              180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241,
              71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_3 (
    .x_in(stage_6_per_out[6]),
    .y_in(stage_6_per_out[7]),
    .x_out(stage_7_per_in[6]),
    .y_out(stage_7_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896,
              180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241,
              71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_4 (
    .x_in(stage_6_per_out[8]),
    .y_in(stage_6_per_out[9]),
    .x_out(stage_7_per_in[8]),
    .y_out(stage_7_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896,
              180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241,
              71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_5 (
    .x_in(stage_6_per_out[10]),
    .y_in(stage_6_per_out[11]),
    .x_out(stage_7_per_in[10]),
    .y_out(stage_7_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896,
              180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241,
              71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_6 (
    .x_in(stage_6_per_out[12]),
    .y_in(stage_6_per_out[13]),
    .x_out(stage_7_per_in[12]),
    .y_out(stage_7_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896,
              180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241,
              71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_7 (
    .x_in(stage_6_per_out[14]),
    .y_in(stage_6_per_out[15]),
    .x_out(stage_7_per_in[14]),
    .y_out(stage_7_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896,
              180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241,
              71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_8 (
    .x_in(stage_6_per_out[16]),
    .y_in(stage_6_per_out[17]),
    .x_out(stage_7_per_in[16]),
    .y_out(stage_7_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896,
              180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241,
              71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_9 (
    .x_in(stage_6_per_out[18]),
    .y_in(stage_6_per_out[19]),
    .x_out(stage_7_per_in[18]),
    .y_out(stage_7_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896,
              180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241,
              71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_10 (
    .x_in(stage_6_per_out[20]),
    .y_in(stage_6_per_out[21]),
    .x_out(stage_7_per_in[20]),
    .y_out(stage_7_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896,
              180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241,
              71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_11 (
    .x_in(stage_6_per_out[22]),
    .y_in(stage_6_per_out[23]),
    .x_out(stage_7_per_in[22]),
    .y_out(stage_7_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896,
              180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241,
              71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_12 (
    .x_in(stage_6_per_out[24]),
    .y_in(stage_6_per_out[25]),
    .x_out(stage_7_per_in[24]),
    .y_out(stage_7_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896,
              180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241,
              71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_13 (
    .x_in(stage_6_per_out[26]),
    .y_in(stage_6_per_out[27]),
    .x_out(stage_7_per_in[26]),
    .y_out(stage_7_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896,
              180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241,
              71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_14 (
    .x_in(stage_6_per_out[28]),
    .y_in(stage_6_per_out[29]),
    .x_out(stage_7_per_in[28]),
    .y_out(stage_7_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896, 96332896,
              180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988, 180609988,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261, 130838261,
              90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588, 90670588,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241, 128108241,
              71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504, 71274504}))
  stage_7_butterfly_15 (
    .x_in(stage_6_per_out[30]),
    .y_in(stage_6_per_out[31]),
    .x_out(stage_7_per_in[30]),
    .y_out(stage_7_per_in[31]),
    .clk(clk),
    .rst(rst)
  );





  // TODO(Yang): stage 7 -> stage 8 permutation
  // FIXME: ignore butterfly units for now.
  stage_7_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_7_8_per (
    .inData_0(stage_7_per_in[0]),
    .inData_1(stage_7_per_in[1]),
    .inData_2(stage_7_per_in[2]),
    .inData_3(stage_7_per_in[3]),
    .inData_4(stage_7_per_in[4]),
    .inData_5(stage_7_per_in[5]),
    .inData_6(stage_7_per_in[6]),
    .inData_7(stage_7_per_in[7]),
    .inData_8(stage_7_per_in[8]),
    .inData_9(stage_7_per_in[9]),
    .inData_10(stage_7_per_in[10]),
    .inData_11(stage_7_per_in[11]),
    .inData_12(stage_7_per_in[12]),
    .inData_13(stage_7_per_in[13]),
    .inData_14(stage_7_per_in[14]),
    .inData_15(stage_7_per_in[15]),
    .inData_16(stage_7_per_in[16]),
    .inData_17(stage_7_per_in[17]),
    .inData_18(stage_7_per_in[18]),
    .inData_19(stage_7_per_in[19]),
    .inData_20(stage_7_per_in[20]),
    .inData_21(stage_7_per_in[21]),
    .inData_22(stage_7_per_in[22]),
    .inData_23(stage_7_per_in[23]),
    .inData_24(stage_7_per_in[24]),
    .inData_25(stage_7_per_in[25]),
    .inData_26(stage_7_per_in[26]),
    .inData_27(stage_7_per_in[27]),
    .inData_28(stage_7_per_in[28]),
    .inData_29(stage_7_per_in[29]),
    .inData_30(stage_7_per_in[30]),
    .inData_31(stage_7_per_in[31]),
    .outData_0(stage_7_per_out[0]),
    .outData_1(stage_7_per_out[1]),
    .outData_2(stage_7_per_out[2]),
    .outData_3(stage_7_per_out[3]),
    .outData_4(stage_7_per_out[4]),
    .outData_5(stage_7_per_out[5]),
    .outData_6(stage_7_per_out[6]),
    .outData_7(stage_7_per_out[7]),
    .outData_8(stage_7_per_out[8]),
    .outData_9(stage_7_per_out[9]),
    .outData_10(stage_7_per_out[10]),
    .outData_11(stage_7_per_out[11]),
    .outData_12(stage_7_per_out[12]),
    .outData_13(stage_7_per_out[13]),
    .outData_14(stage_7_per_out[14]),
    .outData_15(stage_7_per_out[15]),
    .outData_16(stage_7_per_out[16]),
    .outData_17(stage_7_per_out[17]),
    .outData_18(stage_7_per_out[18]),
    .outData_19(stage_7_per_out[19]),
    .outData_20(stage_7_per_out[20]),
    .outData_21(stage_7_per_out[21]),
    .outData_22(stage_7_per_out[22]),
    .outData_23(stage_7_per_out[23]),
    .outData_24(stage_7_per_out[24]),
    .outData_25(stage_7_per_out[25]),
    .outData_26(stage_7_per_out[26]),
    .outData_27(stage_7_per_out[27]),
    .outData_28(stage_7_per_out[28]),
    .outData_29(stage_7_per_out[29]),
    .outData_30(stage_7_per_out[30]),
    .outData_31(stage_7_per_out[31]),
    .in_start(in_start[7]),
    .out_start(out_start[7]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 8 32 butterfly units
  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_0 (
    .x_in(stage_7_per_out[0]),
    .y_in(stage_7_per_out[1]),
    .x_out(stage_8_per_in[0]),
    .y_out(stage_8_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_1 (
    .x_in(stage_7_per_out[2]),
    .y_in(stage_7_per_out[3]),
    .x_out(stage_8_per_in[2]),
    .y_out(stage_8_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_2 (
    .x_in(stage_7_per_out[4]),
    .y_in(stage_7_per_out[5]),
    .x_out(stage_8_per_in[4]),
    .y_out(stage_8_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_3 (
    .x_in(stage_7_per_out[6]),
    .y_in(stage_7_per_out[7]),
    .x_out(stage_8_per_in[6]),
    .y_out(stage_8_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_4 (
    .x_in(stage_7_per_out[8]),
    .y_in(stage_7_per_out[9]),
    .x_out(stage_8_per_in[8]),
    .y_out(stage_8_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_5 (
    .x_in(stage_7_per_out[10]),
    .y_in(stage_7_per_out[11]),
    .x_out(stage_8_per_in[10]),
    .y_out(stage_8_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_6 (
    .x_in(stage_7_per_out[12]),
    .y_in(stage_7_per_out[13]),
    .x_out(stage_8_per_in[12]),
    .y_out(stage_8_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_7 (
    .x_in(stage_7_per_out[14]),
    .y_in(stage_7_per_out[15]),
    .x_out(stage_8_per_in[14]),
    .y_out(stage_8_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_8 (
    .x_in(stage_7_per_out[16]),
    .y_in(stage_7_per_out[17]),
    .x_out(stage_8_per_in[16]),
    .y_out(stage_8_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_9 (
    .x_in(stage_7_per_out[18]),
    .y_in(stage_7_per_out[19]),
    .x_out(stage_8_per_in[18]),
    .y_out(stage_8_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_10 (
    .x_in(stage_7_per_out[20]),
    .y_in(stage_7_per_out[21]),
    .x_out(stage_8_per_in[20]),
    .y_out(stage_8_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_11 (
    .x_in(stage_7_per_out[22]),
    .y_in(stage_7_per_out[23]),
    .x_out(stage_8_per_in[22]),
    .y_out(stage_8_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_12 (
    .x_in(stage_7_per_out[24]),
    .y_in(stage_7_per_out[25]),
    .x_out(stage_8_per_in[24]),
    .y_out(stage_8_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_13 (
    .x_in(stage_7_per_out[26]),
    .y_in(stage_7_per_out[27]),
    .x_out(stage_8_per_in[26]),
    .y_out(stage_8_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_14 (
    .x_in(stage_7_per_out[28]),
    .y_in(stage_7_per_out[29]),
    .x_out(stage_8_per_in[28]),
    .y_out(stage_8_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460, 18186460,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205,
              93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205, 93509205}))
  stage_8_butterfly_15 (
    .x_in(stage_7_per_out[30]),
    .y_in(stage_7_per_out[31]),
    .x_out(stage_8_per_in[30]),
    .y_out(stage_8_per_in[31]),
    .clk(clk),
    .rst(rst)
  );





  // TODO(Yang): stage 8 -> stage 9 permutation
  // FIXME: ignore butterfly units for now.
  stage_8_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_8_9_per (
    .inData_0(stage_8_per_in[0]),
    .inData_1(stage_8_per_in[1]),
    .inData_2(stage_8_per_in[2]),
    .inData_3(stage_8_per_in[3]),
    .inData_4(stage_8_per_in[4]),
    .inData_5(stage_8_per_in[5]),
    .inData_6(stage_8_per_in[6]),
    .inData_7(stage_8_per_in[7]),
    .inData_8(stage_8_per_in[8]),
    .inData_9(stage_8_per_in[9]),
    .inData_10(stage_8_per_in[10]),
    .inData_11(stage_8_per_in[11]),
    .inData_12(stage_8_per_in[12]),
    .inData_13(stage_8_per_in[13]),
    .inData_14(stage_8_per_in[14]),
    .inData_15(stage_8_per_in[15]),
    .inData_16(stage_8_per_in[16]),
    .inData_17(stage_8_per_in[17]),
    .inData_18(stage_8_per_in[18]),
    .inData_19(stage_8_per_in[19]),
    .inData_20(stage_8_per_in[20]),
    .inData_21(stage_8_per_in[21]),
    .inData_22(stage_8_per_in[22]),
    .inData_23(stage_8_per_in[23]),
    .inData_24(stage_8_per_in[24]),
    .inData_25(stage_8_per_in[25]),
    .inData_26(stage_8_per_in[26]),
    .inData_27(stage_8_per_in[27]),
    .inData_28(stage_8_per_in[28]),
    .inData_29(stage_8_per_in[29]),
    .inData_30(stage_8_per_in[30]),
    .inData_31(stage_8_per_in[31]),
    .outData_0(stage_8_per_out[0]),
    .outData_1(stage_8_per_out[1]),
    .outData_2(stage_8_per_out[2]),
    .outData_3(stage_8_per_out[3]),
    .outData_4(stage_8_per_out[4]),
    .outData_5(stage_8_per_out[5]),
    .outData_6(stage_8_per_out[6]),
    .outData_7(stage_8_per_out[7]),
    .outData_8(stage_8_per_out[8]),
    .outData_9(stage_8_per_out[9]),
    .outData_10(stage_8_per_out[10]),
    .outData_11(stage_8_per_out[11]),
    .outData_12(stage_8_per_out[12]),
    .outData_13(stage_8_per_out[13]),
    .outData_14(stage_8_per_out[14]),
    .outData_15(stage_8_per_out[15]),
    .outData_16(stage_8_per_out[16]),
    .outData_17(stage_8_per_out[17]),
    .outData_18(stage_8_per_out[18]),
    .outData_19(stage_8_per_out[19]),
    .outData_20(stage_8_per_out[20]),
    .outData_21(stage_8_per_out[21]),
    .outData_22(stage_8_per_out[22]),
    .outData_23(stage_8_per_out[23]),
    .outData_24(stage_8_per_out[24]),
    .outData_25(stage_8_per_out[25]),
    .outData_26(stage_8_per_out[26]),
    .outData_27(stage_8_per_out[27]),
    .outData_28(stage_8_per_out[28]),
    .outData_29(stage_8_per_out[29]),
    .outData_30(stage_8_per_out[30]),
    .outData_31(stage_8_per_out[31]),
    .in_start(in_start[8]),
    .out_start(out_start[8]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 9 32 butterfly units
  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_0 (
    .x_in(stage_8_per_out[0]),
    .y_in(stage_8_per_out[1]),
    .x_out(stage_9_per_in[0]),
    .y_out(stage_9_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_1 (
    .x_in(stage_8_per_out[2]),
    .y_in(stage_8_per_out[3]),
    .x_out(stage_9_per_in[2]),
    .y_out(stage_9_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_2 (
    .x_in(stage_8_per_out[4]),
    .y_in(stage_8_per_out[5]),
    .x_out(stage_9_per_in[4]),
    .y_out(stage_9_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_3 (
    .x_in(stage_8_per_out[6]),
    .y_in(stage_8_per_out[7]),
    .x_out(stage_9_per_in[6]),
    .y_out(stage_9_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_4 (
    .x_in(stage_8_per_out[8]),
    .y_in(stage_8_per_out[9]),
    .x_out(stage_9_per_in[8]),
    .y_out(stage_9_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_5 (
    .x_in(stage_8_per_out[10]),
    .y_in(stage_8_per_out[11]),
    .x_out(stage_9_per_in[10]),
    .y_out(stage_9_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_6 (
    .x_in(stage_8_per_out[12]),
    .y_in(stage_8_per_out[13]),
    .x_out(stage_9_per_in[12]),
    .y_out(stage_9_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_7 (
    .x_in(stage_8_per_out[14]),
    .y_in(stage_8_per_out[15]),
    .x_out(stage_9_per_in[14]),
    .y_out(stage_9_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_8 (
    .x_in(stage_8_per_out[16]),
    .y_in(stage_8_per_out[17]),
    .x_out(stage_9_per_in[16]),
    .y_out(stage_9_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_9 (
    .x_in(stage_8_per_out[18]),
    .y_in(stage_8_per_out[19]),
    .x_out(stage_9_per_in[18]),
    .y_out(stage_9_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_10 (
    .x_in(stage_8_per_out[20]),
    .y_in(stage_8_per_out[21]),
    .x_out(stage_9_per_in[20]),
    .y_out(stage_9_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_11 (
    .x_in(stage_8_per_out[22]),
    .y_in(stage_8_per_out[23]),
    .x_out(stage_9_per_in[22]),
    .y_out(stage_9_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_12 (
    .x_in(stage_8_per_out[24]),
    .y_in(stage_8_per_out[25]),
    .x_out(stage_9_per_in[24]),
    .y_out(stage_9_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_13 (
    .x_in(stage_8_per_out[26]),
    .y_in(stage_8_per_out[27]),
    .x_out(stage_9_per_in[26]),
    .y_out(stage_9_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_14 (
    .x_in(stage_8_per_out[28]),
    .y_in(stage_8_per_out[29]),
    .x_out(stage_9_per_in[28]),
    .y_out(stage_9_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802}))
  stage_9_butterfly_15 (
    .x_in(stage_8_per_out[30]),
    .y_in(stage_8_per_out[31]),
    .x_out(stage_9_per_in[30]),
    .y_out(stage_9_per_in[31]),
    .clk(clk),
    .rst(rst)
  );


  // TODO(Yang): Update stride
  stage_9_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_9_10_per (
    .inData_0(stage_9_per_in[0]),
    .inData_1(stage_9_per_in[1]),
    .inData_2(stage_9_per_in[2]),
    .inData_3(stage_9_per_in[3]),
    .inData_4(stage_9_per_in[4]),
    .inData_5(stage_9_per_in[5]),
    .inData_6(stage_9_per_in[6]),
    .inData_7(stage_9_per_in[7]),
    .inData_8(stage_9_per_in[8]),
    .inData_9(stage_9_per_in[9]),
    .inData_10(stage_9_per_in[10]),
    .inData_11(stage_9_per_in[11]),
    .inData_12(stage_9_per_in[12]),
    .inData_13(stage_9_per_in[13]),
    .inData_14(stage_9_per_in[14]),
    .inData_15(stage_9_per_in[15]),
    .inData_16(stage_9_per_in[16]),
    .inData_17(stage_9_per_in[17]),
    .inData_18(stage_9_per_in[18]),
    .inData_19(stage_9_per_in[19]),
    .inData_20(stage_9_per_in[20]),
    .inData_21(stage_9_per_in[21]),
    .inData_22(stage_9_per_in[22]),
    .inData_23(stage_9_per_in[23]),
    .inData_24(stage_9_per_in[24]),
    .inData_25(stage_9_per_in[25]),
    .inData_26(stage_9_per_in[26]),
    .inData_27(stage_9_per_in[27]),
    .inData_28(stage_9_per_in[28]),
    .inData_29(stage_9_per_in[29]),
    .inData_30(stage_9_per_in[30]),
    .inData_31(stage_9_per_in[31]),
    .outData_0(stage_9_per_out[0]),
    .outData_1(stage_9_per_out[1]),
    .outData_2(stage_9_per_out[2]),
    .outData_3(stage_9_per_out[3]),
    .outData_4(stage_9_per_out[4]),
    .outData_5(stage_9_per_out[5]),
    .outData_6(stage_9_per_out[6]),
    .outData_7(stage_9_per_out[7]),
    .outData_8(stage_9_per_out[8]),
    .outData_9(stage_9_per_out[9]),
    .outData_10(stage_9_per_out[10]),
    .outData_11(stage_9_per_out[11]),
    .outData_12(stage_9_per_out[12]),
    .outData_13(stage_9_per_out[13]),
    .outData_14(stage_9_per_out[14]),
    .outData_15(stage_9_per_out[15]),
    .outData_16(stage_9_per_out[16]),
    .outData_17(stage_9_per_out[17]),
    .outData_18(stage_9_per_out[18]),
    .outData_19(stage_9_per_out[19]),
    .outData_20(stage_9_per_out[20]),
    .outData_21(stage_9_per_out[21]),
    .outData_22(stage_9_per_out[22]),
    .outData_23(stage_9_per_out[23]),
    .outData_24(stage_9_per_out[24]),
    .outData_25(stage_9_per_out[25]),
    .outData_26(stage_9_per_out[26]),
    .outData_27(stage_9_per_out[27]),
    .outData_28(stage_9_per_out[28]),
    .outData_29(stage_9_per_out[29]),
    .outData_30(stage_9_per_out[30]),
    .outData_31(stage_9_per_out[31]),
    .in_start(in_start[9]),
    .out_start(out_start[9]),
    .clk(clk),
    .rst(rst)
  );

  // TODO(Tian): stage 10 32 butterfly units
  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_0 (
    .x_in(stage_9_per_out[0]),
    .y_in(stage_9_per_out[1]),
    .x_out(outData[0]),
    .y_out(outData[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_1 (
    .x_in(stage_9_per_out[2]),
    .y_in(stage_9_per_out[3]),
    .x_out(outData[2]),
    .y_out(outData[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_2 (
    .x_in(stage_9_per_out[4]),
    .y_in(stage_9_per_out[5]),
    .x_out(outData[4]),
    .y_out(outData[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_3 (
    .x_in(stage_9_per_out[6]),
    .y_in(stage_9_per_out[7]),
    .x_out(outData[6]),
    .y_out(outData[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_4 (
    .x_in(stage_9_per_out[8]),
    .y_in(stage_9_per_out[9]),
    .x_out(outData[8]),
    .y_out(outData[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_5 (
    .x_in(stage_9_per_out[10]),
    .y_in(stage_9_per_out[11]),
    .x_out(outData[10]),
    .y_out(outData[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_6 (
    .x_in(stage_9_per_out[12]),
    .y_in(stage_9_per_out[13]),
    .x_out(outData[12]),
    .y_out(outData[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_7 (
    .x_in(stage_9_per_out[14]),
    .y_in(stage_9_per_out[15]),
    .x_out(outData[14]),
    .y_out(outData[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_8 (
    .x_in(stage_9_per_out[16]),
    .y_in(stage_9_per_out[17]),
    .x_out(outData[16]),
    .y_out(outData[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_9 (
    .x_in(stage_9_per_out[18]),
    .y_in(stage_9_per_out[19]),
    .x_out(outData[18]),
    .y_out(outData[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_10 (
    .x_in(stage_9_per_out[20]),
    .y_in(stage_9_per_out[21]),
    .x_out(outData[20]),
    .y_out(outData[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_11 (
    .x_in(stage_9_per_out[22]),
    .y_in(stage_9_per_out[23]),
    .x_out(outData[22]),
    .y_out(outData[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_12 (
    .x_in(stage_9_per_out[24]),
    .y_in(stage_9_per_out[25]),
    .x_out(outData[24]),
    .y_out(outData[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_13 (
    .x_in(stage_9_per_out[26]),
    .y_in(stage_9_per_out[27]),
    .x_out(outData[26]),
    .y_out(outData[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_14 (
    .x_in(stage_9_per_out[28]),
    .y_in(stage_9_per_out[29]),
    .x_out(outData[28]),
    .y_out(outData[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761,
              75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761, 75074761}))
  stage_10_butterfly_15 (
    .x_in(stage_9_per_out[30]),
    .y_in(stage_9_per_out[31]),
    .x_out(outData[30]),
    .y_out(outData[31]),
    .clk(clk),
    .rst(rst)
  );


endmodule
