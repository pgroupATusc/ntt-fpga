// NTT Accelerator

module NTT_Top #(
    parameter NUM_BITS_PER_INPUT = 32
  ) (
    clk,
    rst,
    ...
  );

endmodule
