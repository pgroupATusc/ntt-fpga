// NTT Accelerator

module NTT_Top #(
    parameter DATA_WIDTH_PER_INPUT = 28,
    parameter INPUT_PER_CYCLE = 32
  ) (
    inData,
    outData,
    in_start,
    out_start,
    clk,
    rst,
  );

  input clk, rst;

  input in_start[10:0];
  output logic out_start[10:0];

  input        [DATA_WIDTH_PER_INPUT-1:0] inData[INPUT_PER_CYCLE-1:0];
  output logic [DATA_WIDTH_PER_INPUT-1:0] outData[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_0_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_0_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_1_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_1_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_2_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_2_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_3_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_3_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_4_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_4_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_5_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_5_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_6_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_6_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_7_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_7_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_8_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_8_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_9_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_9_per_out[INPUT_PER_CYCLE-1:0];

  logic [DATA_WIDTH_PER_INPUT-1:0] stage_10_per_in[INPUT_PER_CYCLE-1:0];
  logic [DATA_WIDTH_PER_INPUT-1:0] stage_10_per_out[INPUT_PER_CYCLE-1:0];

  parameter [8:0] START_CYCLE[12] = {0, 7, 14, 21, 28, 49, 71, 95, 123, 159, 211, 295};

  // TODO(Tian): stage 0 32 butterfly units
  butterfly #(
    .start(START_CYCLE[0]),
    .factors({62736, 138390585, 229351752, 232397550, 248258143, 237695631, 5986200, 76613625,
              141200910, 260020495, 238271990, 251656189, 210432655, 47407140, 139336311, 30182006,
              60410137, 50557363, 227274721, 225306517, 60657405, 63634221, 217306794, 173443464,
              120438379, 126074738, 125625707, 115237475, 154088507, 131255494, 162143577, 75233812,
              168799557, 209093018, 115574858, 85762236, 163194978, 214996992, 4369826, 59403344,
              90751938, 159528330, 24738255, 174916329, 174394830, 39518152, 21511271, 238064453,
              65612009, 221285249, 151945076, 16499278, 26268761, 71341164, 224561048, 81430431,
              42684255, 171732518, 135812431, 202855239, 178512370, 73723002, 96512966, 2615849,
              8259075, 69789389, 86907964, 1371159, 229881708, 114463563, 233570711, 196480564,
              81393489, 219691960, 136863777, 139897823, 184579826, 262334367, 193086087, 199105134,
              66137976, 229237307, 46407972, 49661599, 168246811, 253577157, 9971642, 33454619,
              131575231, 127322073, 215932086, 360580, 114248229, 126370638, 132028761, 85118780,
              104041706, 103557733, 228870065, 215247918, 39123511, 187113601, 173212060, 172102431,
              110271140, 55682893, 130565708, 234938972, 151231163, 256536575, 147718178, 13664359,
              9497918, 123998976, 131123953, 18799530, 10785136, 258162508, 167082925, 242453874,
              146990305, 228964332, 12430538, 197777956, 228578092, 108727234, 263121861, 261712272}))
  stage_0_butterfly_0 (
    .x_in(inData[0]),
    .y_in(inData[1]),
    .x_out(stage_0_per_in[0]),
    .y_out(stage_0_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({1907454, 18568532, 18284087, 173978412, 179300118, 142538555, 3778321, 183539945,
              190023698, 73697328, 215835949, 35857213, 238852009, 53030863, 79816727, 202544817,
              90459251, 148940015, 38780522, 152136534, 188631715, 148753884, 180949546, 107281991,
              93000404, 35553140, 179673158, 220692949, 68711843, 249640388, 48588607, 135453164,
              145932355, 196709411, 25746466, 145101039, 136072729, 252862876, 68336365, 56280600,
              125408694, 194605816, 31768873, 236121751, 234613484, 241597278, 42275209, 254006109,
              18646649, 121142478, 82056103, 267007570, 241285957, 206826789, 195819103, 41756449,
              249490832, 147507351, 22776264, 87928571, 138558999, 240078055, 241947117, 13493318,
              224650429, 229741385, 132709741, 21489734, 75771663, 196341244, 106442355, 187504892,
              118813697, 217792655, 213823426, 247808775, 184231755, 120846747, 222306946, 28244848,
              48524018, 86285917, 6841080, 208868555, 184001594, 182145624, 59811701, 79440456,
              149996455, 48555419, 108455048, 16609890, 9255299, 2353936, 122257237, 59625292,
              70352813, 160793918, 244570986, 1618864, 49444600, 110273227, 48810421, 205236559,
              34248663, 126498799, 35295690, 46583536, 236243144, 136554164, 231200794, 99167958,
              125590824, 57499821, 182424131, 74632878, 135108737, 53524475, 84704450, 167937680,
              176139969, 86892569, 232516826, 167199557, 129357001, 244434992, 17124429, 142049175}))
  stage_0_butterfly_1 (
    .x_in(inData[2]),
    .y_in(inData[3]),
    .x_out(stage_0_per_in[2]),
    .y_out(stage_0_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({127608977, 5473511, 121332251, 266521776, 157389868, 144769477, 3052481, 21572447,
              238966374, 46912433, 154495952, 56987360, 172782070, 26866408, 49806007, 94223513,
              127870778, 213245383, 70554670, 20426733, 249304086, 85422012, 54418504, 66819851,
              229943365, 150130406, 135886727, 181022773, 896607, 169515998, 41484727, 203722503,
              111929529, 132349487, 235715975, 75105065, 41726718, 221059178, 27836602, 2011982,
              264371342, 11959677, 149329993, 129605716, 198700251, 219029055, 228606302, 7229020,
              140808004, 9479322, 25249547, 206462525, 155953488, 27115908, 212109347, 234710989,
              105651651, 36246851, 24888645, 107677384, 95350060, 212385093, 158561039, 194562323,
              190509603, 130771778, 260134415, 49717914, 169809008, 163019788, 236342274, 66144131,
              251686044, 107104549, 130863524, 173951180, 218474935, 107135677, 244025737, 246477773,
              65316150, 44515532, 51724689, 251263130, 179814135, 263884483, 47156256, 185730304,
              122737973, 162829016, 108348559, 14692215, 239606434, 251425486, 183216854, 255690434,
              221042295, 87325743, 267488469, 112251860, 186854087, 211366667, 198490305, 158126231,
              15301013, 86460683, 97252224, 153141493, 24230656, 151221429, 109429555, 229582731,
              104126955, 11703135, 7378856, 100946881, 72034061, 106563970, 140793205, 34699254,
              83950689, 177264548, 254596309, 149344309, 184896958, 225116841, 27247099, 151842442}))
  stage_0_butterfly_2 (
    .x_in(inData[4]),
    .y_in(inData[5]),
    .x_out(stage_0_per_in[4]),
    .y_out(stage_0_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({169184935, 125480909, 106831467, 184791819, 195652857, 5231854, 14448911, 151524267,
              91778054, 81083779, 36311778, 56333048, 32605484, 265950738, 152480704, 179139190,
              129584651, 81873483, 110996066, 186348595, 223960411, 4986407, 45577523, 8297893,
              35630094, 155163691, 68771072, 109371065, 255719214, 208653574, 48342959, 213678319,
              123658638, 112142792, 154830655, 174632895, 202025824, 96892627, 121686109, 258549338,
              210012123, 55192006, 260828874, 194603131, 140340588, 60603436, 245765723, 28116292,
              170942291, 155517338, 125238212, 66449840, 215941659, 260087354, 20537000, 255738903,
              132315280, 90006293, 129408474, 188542273, 102742547, 242826313, 44845193, 78592957,
              180416915, 100132307, 237936557, 5068353, 30247571, 210363951, 122360079, 96374025,
              104447750, 164529221, 5132066, 29805745, 197344625, 202640881, 13810215, 197497401,
              194219704, 256480283, 162923321, 231677557, 32737194, 123317306, 103204044, 230350716,
              188122907, 6725515, 217085295, 69230198, 179717207, 218852619, 92792804, 4491002,
              72945707, 135171113, 143112792, 116647317, 210644544, 9249520, 152283243, 244555167,
              249388588, 128889378, 60682421, 90584256, 181705475, 242671835, 33223660, 47508483,
              107928332, 48777982, 119835732, 179869441, 77051365, 30822536, 150857390, 175007080,
              46671057, 188656071, 122169973, 43714082, 12667818, 56125789, 34847782, 136274746}))
  stage_0_butterfly_3 (
    .x_in(inData[6]),
    .y_in(inData[7]),
    .x_out(stage_0_per_in[6]),
    .y_out(stage_0_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({221849129, 234869713, 151923798, 260851907, 74962493, 226595737, 133797910, 42776728,
              40496733, 206537906, 2862602, 39521553, 229751485, 189986560, 117960054, 194846985,
              173052617, 42053510, 105948718, 15379209, 254027033, 211444110, 20059876, 61891902,
              200934478, 208159538, 26464113, 254332699, 77856633, 242184182, 182951273, 192707093,
              41023501, 234287689, 34644106, 105706660, 61497280, 76639397, 265346073, 152738846,
              230823778, 228971558, 131105010, 37752789, 170978026, 245369685, 44078325, 142898101,
              132556999, 41652472, 47307859, 158858535, 24970434, 95816060, 79305722, 145592959,
              136104512, 82875459, 205576016, 185232992, 61680409, 259733399, 192247464, 204313060,
              143100858, 186545936, 233222120, 260923957, 163860332, 261016176, 134390440, 134614101,
              181610634, 243862110, 153531059, 176789033, 76430728, 112718220, 101462472, 97251575,
              181981633, 50106798, 232770856, 13704349, 98483239, 84901432, 57501675, 222748125,
              207033531, 229222177, 46461494, 109746000, 228091235, 90105969, 24794247, 263215622,
              8255313, 266284483, 238036964, 69414413, 200339141, 148796874, 59294895, 42275800,
              170921357, 135646873, 118725672, 207530553, 158126817, 148098547, 110117913, 69218942,
              38773847, 166068773, 167554606, 53167918, 171975768, 244602309, 84361140, 150154963,
              247783732, 99177320, 188917923, 110104975, 69921988, 255918779, 78030852, 57302073}))
  stage_0_butterfly_4 (
    .x_in(inData[8]),
    .y_in(inData[9]),
    .x_out(stage_0_per_in[8]),
    .y_out(stage_0_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({172988180, 250606181, 185050869, 29470818, 67529023, 149138685, 104771116, 54233307,
              41146808, 240784947, 129899073, 132129988, 88521257, 158533760, 225676034, 248896168,
              90342181, 212167090, 243834156, 27029386, 203523838, 228871862, 156432226, 26659480,
              234989972, 205287356, 116017893, 176832880, 49058740, 61691447, 247983171, 258883039,
              51002920, 109505067, 255155441, 21131779, 18305869, 35559942, 12986586, 66715025,
              67916891, 240649845, 231410375, 229784592, 225077819, 62782868, 215954984, 115679885,
              72252210, 159471860, 112561771, 153682120, 143573525, 235388028, 227071465, 59375296,
              81013691, 230143339, 119190794, 186483628, 243451530, 143816111, 60134449, 72475326,
              124282928, 12651571, 131237870, 157068444, 198223, 244905743, 249630983, 54358169,
              18803294, 175334429, 201861189, 260001724, 253464518, 59370938, 107586283, 209246609,
              129798040, 58677377, 186098576, 113781795, 185094855, 249212399, 239753050, 77840672,
              265171130, 225914175, 158309971, 179365619, 160882583, 38752877, 192193505, 7116217,
              62374498, 236327891, 219418748, 263718984, 154596247, 157430256, 32372991, 158711864,
              168351315, 233906629, 33508832, 74385386, 263412265, 20877990, 106358666, 198306293,
              118482368, 220394580, 157437159, 152365066, 248278309, 198378776, 38642987, 245615084,
              26045295, 265616179, 248241093, 192872385, 36987199, 260374016, 144111858, 72549374}))
  stage_0_butterfly_5 (
    .x_in(inData[10]),
    .y_in(inData[11]),
    .x_out(stage_0_per_in[10]),
    .y_out(stage_0_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({163149532, 5740730, 94277220, 167586303, 144055138, 218879515, 228780544, 112058009,
              120515996, 116970950, 12984872, 63216411, 55158081, 104949331, 157537739, 132200486,
              69936597, 42733910, 63986967, 83981669, 215111514, 197423642, 171719097, 12855237,
              44459414, 128505750, 184499901, 171842488, 150205042, 96976591, 152039665, 96526884,
              227615757, 151704879, 110912131, 27233477, 246680455, 154775650, 182209928, 264329231,
              6265971, 109376139, 223045283, 82632268, 110327668, 162925843, 235787722, 21764948,
              50475029, 31551002, 36214289, 144184457, 259992880, 13842453, 14462331, 235284227,
              65760618, 181725973, 54697818, 83931467, 161245819, 132907662, 259993096, 97581367,
              87220148, 63656435, 68196879, 136382259, 39654333, 230967163, 199075664, 2029098,
              81207363, 149477651, 76114224, 254244111, 7447708, 185120393, 120912967, 102116116,
              81762412, 234954565, 106463701, 227944808, 120134099, 46729148, 227158983, 89270439,
              252263799, 24734017, 170302338, 213642756, 71887650, 108647642, 228212013, 212003953,
              122977291, 150283834, 144673958, 61250374, 519479, 67046513, 123713876, 2557700,
              59384117, 136400329, 178886927, 170944566, 118024210, 28935497, 199074208, 202918045,
              110162160, 99410963, 112635657, 206482017, 79702710, 134843781, 213908547, 235546264,
              17550542, 108704486, 93347053, 117771098, 132702632, 41112252, 17823318, 220194496}))
  stage_0_butterfly_6 (
    .x_in(inData[12]),
    .y_in(inData[13]),
    .x_out(stage_0_per_in[12]),
    .y_out(stage_0_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({196855462, 179625763, 128643267, 148827249, 205246482, 21458183, 224318864, 1696019,
              131370540, 88419162, 131972043, 58280814, 68756958, 81930, 205821112, 131559431,
              97670877, 70436067, 34174616, 192680584, 39872790, 184608754, 265191298, 13429213,
              162528302, 39140268, 51441041, 39919904, 170882254, 211152508, 171967455, 115525972,
              138161289, 234322267, 3764785, 213843114, 200939178, 111908324, 113870289, 17233293,
              234685655, 243297654, 66804322, 262250139, 210089549, 78892295, 218637579, 173572777,
              258291717, 246940389, 92763586, 162490819, 105582618, 192516565, 222708254, 82054424,
              176214933, 194815301, 234300746, 108661782, 57174663, 147106083, 259999423, 157468594,
              7092568, 88702124, 79425600, 97492082, 37710032, 59212137, 39822794, 234121810,
              267102876, 159725962, 242814722, 156378126, 145439741, 145355888, 108148659, 185671812,
              162088178, 35430665, 194119116, 164207528, 193601964, 27694231, 28536923, 78696193,
              37647978, 180249606, 57720967, 204398753, 221029739, 70151518, 195919352, 99516991,
              7571096, 21742303, 227038693, 116801865, 23520122, 212770879, 28811566, 230635721,
              225275209, 106511467, 161625502, 15750398, 164281505, 171241703, 122116963, 202001175,
              156290837, 231268416, 185167965, 130387641, 1058331, 187415781, 117333915, 37225330,
              173307030, 138920976, 193454786, 18191490, 100165037, 179287997, 83862241, 159562860}))
  stage_0_butterfly_7 (
    .x_in(inData[14]),
    .y_in(inData[15]),
    .x_out(stage_0_per_in[14]),
    .y_out(stage_0_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({58836748, 106056773, 155464901, 48491280, 229152485, 208950205, 255568559, 6668530,
              37016200, 239404299, 757759, 24825329, 30197592, 263982663, 130707805, 185532067,
              198671577, 240039943, 137536510, 136783171, 155288254, 57437223, 237348335, 211688613,
              75750547, 100943177, 141768337, 209177739, 151080366, 4470762, 223003866, 41306715,
              24825033, 136599943, 176371562, 24132582, 244557461, 18792168, 217608608, 146607869,
              164519211, 179831843, 183965087, 111072250, 98922830, 212470099, 267382061, 208828758,
              53079368, 7369182, 49387461, 171197489, 244197291, 144151142, 64306041, 168472713,
              144216104, 116861206, 30614038, 58714599, 189539329, 134997518, 119248989, 206941931,
              215423485, 50402804, 42144250, 183351284, 99315902, 45294283, 221060093, 44427932,
              196350608, 124269051, 208391395, 233581580, 206880652, 168938760, 31181321, 130959181,
              187622314, 159543175, 169601951, 215737735, 15282852, 25904197, 131574531, 84557377,
              191761352, 223537938, 68378584, 165004785, 57198083, 151696189, 146240700, 10658994,
              228922625, 106146355, 209673396, 7620297, 245682235, 213752765, 51270543, 223629100,
              149687609, 3104477, 233335722, 165252821, 135933105, 204917473, 49462279, 38635824,
              90978272, 152734723, 8257788, 264133989, 14827383, 89201641, 212712674, 76772605,
              264868967, 10598408, 239144038, 141503129, 222406475, 164702238, 126093548, 166754761}))
  stage_0_butterfly_8 (
    .x_in(inData[16]),
    .y_in(inData[17]),
    .x_out(stage_0_per_in[16]),
    .y_out(stage_0_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({214715735, 58136368, 235762007, 268021045, 196177971, 201838233, 205271224, 155885829,
              240473245, 170979076, 211663060, 194935198, 180175431, 63162591, 109711544, 103408097,
              238901161, 83840449, 16804445, 216659963, 199052238, 248573392, 95429977, 190439637,
              56018142, 225546029, 174653765, 155010430, 99860276, 15349425, 104275953, 239742054,
              142361011, 177927774, 214327170, 66663233, 182231238, 201356021, 39463122, 179809501,
              223844182, 113458040, 260789685, 201979579, 250127237, 6044206, 130842873, 206641346,
              231138525, 184067420, 32828004, 127364429, 247510253, 70489814, 60661841, 14129846,
              150440065, 136415646, 155312683, 53126633, 158154241, 204076371, 149391390, 134053105,
              71354371, 118651137, 230428614, 111920700, 151814684, 98566622, 106186088, 132259857,
              14667453, 125694138, 69502239, 231794807, 243146642, 107070533, 215911494, 157805049,
              58468223, 250060684, 262471786, 227465231, 94554508, 90061976, 101824639, 27951846,
              250276575, 47826324, 131432446, 168435324, 215943874, 226717406, 225035437, 246208472,
              158081289, 61116726, 192333550, 235669313, 101905032, 120964758, 8718982, 52189384,
              51995938, 136046821, 15958207, 40354434, 82860468, 165567634, 71806036, 131200140,
              264370556, 169435715, 232696276, 203745198, 235758123, 24603905, 60363770, 13532798,
              103662145, 123887389, 262883371, 237430063, 183106668, 55517835, 41823032, 23085612}))
  stage_0_butterfly_9 (
    .x_in(inData[18]),
    .y_in(inData[19]),
    .x_out(stage_0_per_in[18]),
    .y_out(stage_0_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({102340758, 104423755, 160425732, 68227492, 129084525, 189611269, 189138314, 73017801,
              183756330, 21594518, 139937724, 9880764, 57131388, 225369254, 157541500, 156474406,
              39614141, 264479828, 225441652, 127467506, 256641060, 16955107, 97602587, 169350110,
              36695937, 183488163, 190364932, 32128041, 74424009, 179315380, 43784819, 60805498,
              173921335, 27503451, 244546293, 52676293, 233895150, 171672871, 67840088, 83253386,
              237799186, 122367942, 164954582, 172273878, 252406953, 104310584, 238836046, 223368694,
              21531862, 33019077, 62948694, 83749497, 40943954, 156153949, 110250618, 56381879,
              20254495, 241508336, 109921777, 138905259, 21576501, 205242093, 123166625, 221722750,
              164861991, 195906424, 67538787, 107691461, 70654895, 9245191, 152866160, 51218933,
              101813716, 184151583, 194581013, 137830340, 152512971, 236547476, 206403026, 232729335,
              42011142, 67287217, 250005524, 195074984, 166506519, 129666909, 224168732, 4952604,
              251811489, 172140914, 138660240, 16462324, 25877458, 176366269, 14626898, 55752506,
              181180691, 188909348, 135180292, 253757449, 94423638, 230339059, 164438829, 73689066,
              147769827, 16063721, 38284008, 169231043, 115791483, 54766528, 195002054, 205614247,
              242430855, 241821884, 195655909, 95072757, 164243806, 254310437, 5958674, 264371786,
              124253615, 210853880, 192960909, 230124651, 157152581, 221585216, 219422045, 207505578}))
  stage_0_butterfly_10 (
    .x_in(inData[20]),
    .y_in(inData[21]),
    .x_out(stage_0_per_in[20]),
    .y_out(stage_0_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({143786732, 136664320, 75642576, 135770551, 149881682, 224508026, 257328955, 92074820,
              107655283, 92366490, 234828316, 203810197, 81142751, 78969227, 174801883, 91588944,
              159482341, 139852785, 112432362, 62704870, 134571988, 204252016, 114891230, 236052416,
              110693156, 106354792, 122092755, 259685293, 185341670, 168672066, 59653503, 171138130,
              15577361, 81860583, 229528882, 134876482, 180088236, 111274912, 76662541, 55730854,
              183904649, 133008104, 159491283, 152468473, 195538071, 99112512, 204649844, 26767263,
              256986339, 99821278, 87947919, 92092447, 255534095, 34336755, 6777444, 168849030,
              45130170, 216240230, 48856734, 87141435, 129933587, 69177824, 15637687, 96021565,
              88993292, 181033780, 81695275, 201880574, 30549918, 59669292, 261699407, 160584715,
              39931217, 245310720, 237626776, 2176252, 88157673, 138198441, 190689455, 248617642,
              259337446, 106129670, 16392555, 180394230, 51111850, 101060936, 163665671, 229121016,
              256691758, 105408561, 218881712, 171482266, 107087275, 129184142, 72197923, 183002860,
              231263484, 194876189, 243770087, 40301047, 264251329, 74816213, 48869357, 73137377,
              103488513, 71660202, 202431138, 28921814, 172857441, 185723977, 99585718, 152308098,
              11569899, 205958875, 170722015, 30940476, 164573784, 83294274, 63257907, 154688443,
              158386056, 242290819, 152845826, 144681042, 65110284, 163860385, 214283023, 234273255}))
  stage_0_butterfly_11 (
    .x_in(inData[22]),
    .y_in(inData[23]),
    .x_out(stage_0_per_in[22]),
    .y_out(stage_0_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({98227373, 63355713, 26796856, 198563101, 29023980, 224551623, 166961287, 244373783,
              161075491, 89303497, 162545174, 198839540, 23882789, 59001681, 26873848, 227953669,
              22558678, 265709143, 264550106, 135413478, 122229583, 58605619, 157511077, 118174461,
              74718485, 6291440, 246646236, 36389566, 104073065, 146899744, 103787038, 213475348,
              128356119, 260400385, 29220817, 245230909, 38864951, 209546662, 118901157, 170534402,
              178784227, 184276602, 13711872, 158032303, 173580392, 234070704, 156914260, 190758660,
              207607705, 102903513, 198369788, 115048608, 119226838, 224670583, 240151518, 203514552,
              155144532, 45907501, 95898316, 62285640, 208507211, 56939589, 148505031, 150485586,
              239045807, 65941195, 172925747, 43314683, 154170583, 93988508, 97938637, 265006255,
              84715346, 68363059, 34838492, 197478524, 2673613, 19830371, 122693765, 110482921,
              214985679, 85558096, 61883556, 67824335, 113130535, 141580746, 65736109, 135142897,
              22397447, 98503463, 231672458, 174146267, 201302943, 160170338, 110197348, 183449518,
              220005950, 79129285, 32796042, 96257044, 241396543, 124727876, 207300441, 218509565,
              174624298, 291007, 240095534, 227652594, 77968856, 255492938, 89434836, 148811231,
              68807490, 237882452, 49704806, 74916156, 209917670, 8009648, 221163181, 251093184,
              217428510, 127215407, 117652871, 140577689, 193565392, 83000954, 86822274, 34079608}))
  stage_0_butterfly_12 (
    .x_in(inData[24]),
    .y_in(inData[25]),
    .x_out(stage_0_per_in[24]),
    .y_out(stage_0_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({150057464, 101375441, 192174913, 95052731, 23448732, 83959851, 205181101, 112531453,
              101070463, 142276463, 200114, 85927424, 63098068, 228944741, 187534499, 215784466,
              209153008, 147276523, 188446087, 167238213, 144072998, 175168807, 77858155, 230885966,
              247373572, 22914950, 78932104, 196216182, 210239547, 137992276, 268045200, 19847969,
              122550241, 130985550, 54047719, 249112263, 183262830, 198284911, 86866558, 215285662,
              71749872, 175012394, 245038497, 178662179, 180231688, 152315952, 2963416, 154802450,
              134429657, 118213444, 113738086, 40802701, 42021864, 4622329, 247726047, 201888697,
              12808954, 153503748, 77729422, 113731328, 128052742, 225486456, 212184418, 68532350,
              126302082, 107657151, 108404040, 200590842, 6014167, 216371534, 160990548, 255059903,
              78210348, 136530068, 192227833, 214972665, 252922274, 35417568, 162344188, 202258967,
              182834104, 105733032, 225219172, 23130727, 201087126, 7430278, 239353906, 246714101,
              31027015, 41771488, 127805784, 208345113, 42785182, 30147565, 259103093, 23277706,
              33967221, 258487225, 263029881, 117177606, 48087349, 32948426, 169234006, 57795922,
              181325168, 177554441, 23443169, 161226237, 139454911, 68094050, 77508945, 82689315,
              212592244, 149425076, 240905155, 195813478, 170346650, 117454680, 51005918, 44226281,
              108779799, 82939526, 83563004, 208881897, 89733363, 117458270, 193603540, 171515704}))
  stage_0_butterfly_13 (
    .x_in(inData[26]),
    .y_in(inData[27]),
    .x_out(stage_0_per_in[26]),
    .y_out(stage_0_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({39962754, 173776705, 83421235, 37560959, 256558777, 130521421, 14751178, 218305863,
              229530055, 149796825, 110070131, 37761143, 76671502, 167654012, 71449616, 25592978,
              260875356, 69963660, 160647513, 177400482, 10696564, 242086614, 217600940, 125945553,
              25642441, 154162735, 260649789, 88343680, 109410131, 163943008, 175074447, 41373747,
              53554883, 96784305, 114016424, 27425418, 103692636, 178609958, 213474870, 99694466,
              116165973, 183166375, 179512630, 239054686, 51440403, 264712232, 188754097, 137079211,
              266139878, 42583023, 51323950, 177007616, 216328989, 237453043, 247259809, 237567768,
              173030765, 68847542, 65690883, 200029177, 114527376, 245228415, 222486214, 257632808,
              184347612, 17252496, 116203844, 236356015, 32820960, 20606850, 33884144, 148722321,
              176100532, 97520605, 5695672, 50703780, 165433235, 151289170, 140975706, 113484891,
              163077087, 111517965, 135684892, 26760307, 89278624, 41328094, 101029591, 11562888,
              256453055, 140190159, 106059530, 224658359, 149191288, 82596723, 23651884, 130055322,
              197994960, 268107376, 119415929, 625780, 138451058, 92713113, 141473040, 215495577,
              138996529, 217198560, 26132679, 89497967, 151037716, 44239577, 12259140, 211488291,
              49876629, 163847221, 145011041, 216947907, 220416699, 13484173, 148939130, 246176063,
              1235353, 48025256, 135766208, 42743336, 183088464, 95081716, 212842425, 76694868}))
  stage_0_butterfly_14 (
    .x_in(inData[28]),
    .y_in(inData[29]),
    .x_out(stage_0_per_in[28]),
    .y_out(stage_0_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[0]),
    .factors({93261610, 99627052, 141812320, 17746678, 172289773, 36284828, 197944250, 145182880,
              254832984, 193094875, 27854761, 235736575, 258988459, 106508361, 5510115, 228413454,
              108081889, 178085825, 126711917, 10710243, 255307412, 67348921, 59249925, 216347827,
              240106988, 120761900, 86311355, 45256937, 231600531, 247160596, 103407625, 32751373,
              159792872, 150225643, 266701659, 143680187, 94389433, 241625831, 212384234, 192995301,
              126904432, 139998882, 55935675, 168382927, 211721600, 267141235, 52557249, 139421138,
              53728083, 249903585, 205947916, 209077448, 91288416, 259081121, 50951254, 103000049,
              78692480, 134859556, 154254400, 3595020, 122077322, 163361339, 56197115, 99532395,
              16344528, 26620819, 81573675, 134045502, 88484653, 32461064, 117319528, 83014713,
              187760701, 98179318, 95352696, 91252917, 132336250, 213289884, 21476942, 250977019,
              203097121, 226850270, 80678005, 17172477, 158896498, 68554215, 21249308, 101673356,
              185758640, 216246538, 258599303, 161740894, 215878737, 124135460, 114109699, 90052819,
              39817818, 74278900, 44100750, 17691838, 36500136, 97283065, 23918814, 266251087,
              34527937, 118163582, 258759731, 213947035, 116889475, 159360601, 95430596, 134709760,
              138868638, 192889387, 11447146, 1741916, 196733737, 65815578, 103235635, 45566469,
              251183310, 58580381, 180375437, 107220558, 167274958, 239548624, 58071796, 127926589}))
  stage_0_butterfly_15 (
    .x_in(inData[30]),
    .y_in(inData[31]),
    .x_out(stage_0_per_in[30]),
    .y_out(stage_0_per_in[31]),
    .clk(clk),
    .rst(rst)
  );




  // TODO(Yang): stage 0 -> stage 1 permutation
  // FIXME: ignore butterfly units for now.
  stage_0_permutation #(
    .DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    .INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_0_1_per (
    .inData_0(stage_0_per_in[0]),
    .inData_1(stage_0_per_in[1]),
    .inData_2(stage_0_per_in[2]),
    .inData_3(stage_0_per_in[3]),
    .inData_4(stage_0_per_in[4]),
    .inData_5(stage_0_per_in[5]),
    .inData_6(stage_0_per_in[6]),
    .inData_7(stage_0_per_in[7]),
    .inData_8(stage_0_per_in[8]),
    .inData_9(stage_0_per_in[9]),
    .inData_10(stage_0_per_in[10]),
    .inData_11(stage_0_per_in[11]),
    .inData_12(stage_0_per_in[12]),
    .inData_13(stage_0_per_in[13]),
    .inData_14(stage_0_per_in[14]),
    .inData_15(stage_0_per_in[15]),
    .inData_16(stage_0_per_in[16]),
    .inData_17(stage_0_per_in[17]),
    .inData_18(stage_0_per_in[18]),
    .inData_19(stage_0_per_in[19]),
    .inData_20(stage_0_per_in[20]),
    .inData_21(stage_0_per_in[21]),
    .inData_22(stage_0_per_in[22]),
    .inData_23(stage_0_per_in[23]),
    .inData_24(stage_0_per_in[24]),
    .inData_25(stage_0_per_in[25]),
    .inData_26(stage_0_per_in[26]),
    .inData_27(stage_0_per_in[27]),
    .inData_28(stage_0_per_in[28]),
    .inData_29(stage_0_per_in[29]),
    .inData_30(stage_0_per_in[30]),
    .inData_31(stage_0_per_in[31]),
    .outData_0(stage_0_per_out[0]),
    .outData_1(stage_0_per_out[1]),
    .outData_2(stage_0_per_out[2]),
    .outData_3(stage_0_per_out[3]),
    .outData_4(stage_0_per_out[4]),
    .outData_5(stage_0_per_out[5]),
    .outData_6(stage_0_per_out[6]),
    .outData_7(stage_0_per_out[7]),
    .outData_8(stage_0_per_out[8]),
    .outData_9(stage_0_per_out[9]),
    .outData_10(stage_0_per_out[10]),
    .outData_11(stage_0_per_out[11]),
    .outData_12(stage_0_per_out[12]),
    .outData_13(stage_0_per_out[13]),
    .outData_14(stage_0_per_out[14]),
    .outData_15(stage_0_per_out[15]),
    .outData_16(stage_0_per_out[16]),
    .outData_17(stage_0_per_out[17]),
    .outData_18(stage_0_per_out[18]),
    .outData_19(stage_0_per_out[19]),
    .outData_20(stage_0_per_out[20]),
    .outData_21(stage_0_per_out[21]),
    .outData_22(stage_0_per_out[22]),
    .outData_23(stage_0_per_out[23]),
    .outData_24(stage_0_per_out[24]),
    .outData_25(stage_0_per_out[25]),
    .outData_26(stage_0_per_out[26]),
    .outData_27(stage_0_per_out[27]),
    .outData_28(stage_0_per_out[28]),
    .outData_29(stage_0_per_out[29]),
    .outData_30(stage_0_per_out[30]),
    .outData_31(stage_0_per_out[31]),
    .in_start(in_start[0]),
    .out_start(out_start[0]),
    .clk(clk),
    .rst(rst)
  );

  // TODO(Tian): stage 1 32 butterfly units
  butterfly #(
    .start(START_CYCLE[1]),
    .factors({178626802, 22329094, 36426289, 150629496, 226568978, 146360154, 228368554, 175887545,
              142863934, 70370832, 98446051, 171269635, 100723721, 124927121, 195462811, 236561162,
              25937392, 43396787, 48496256, 213843220, 26964940, 37292607, 236960516, 91188581,
              49890248, 52859373, 58870518, 108521058, 57740084, 41918325, 148535761, 67911621,
              238700391, 224183590, 170998790, 104486975, 81363847, 129161289, 54281363, 100791881,
              185850221, 67400723, 153913781, 247062782, 35411505, 48447796, 90710559, 211284483,
              135389110, 260125445, 26451456, 46126435, 34884345, 199208092, 189299702, 222236846,
              212020732, 157341419, 50385541, 31157387, 214331009, 246555646, 46629005, 38115064,
              200295213, 72618725, 6208689, 145706676, 154135831, 222840723, 99461488, 106939991,
              156023579, 116859647, 47430573, 264758616, 139714595, 184120139, 143466178, 17337072,
              214078274, 38429557, 118216948, 195763450, 264282458, 253615348, 173116375, 3677235,
              197485473, 236609676, 9453674, 126894636, 167134668, 19066791, 157049837, 66528431,
              245518247, 53251080, 43737855, 179997990, 195063937, 41015351, 264289232, 81431484,
              205675156, 64307891, 54092187, 204816575, 251274354, 167135704, 198072981, 91524025,
              44349942, 254723792, 100770703, 75117738, 120419308, 147133292, 224620084, 141917139,
              75240990, 4884476, 267404879, 254692251, 143647295, 124656108, 133881133, 45684920}))
  stage_1_butterfly_0 (
    .x_in(stage_0_per_out[0]),
    .y_in(stage_0_per_out[1]),
    .x_out(stage_1_per_in[0]),
    .y_out(stage_1_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({178626802, 22329094, 36426289, 150629496, 226568978, 146360154, 228368554, 175887545,
              142863934, 70370832, 98446051, 171269635, 100723721, 124927121, 195462811, 236561162,
              25937392, 43396787, 48496256, 213843220, 26964940, 37292607, 236960516, 91188581,
              49890248, 52859373, 58870518, 108521058, 57740084, 41918325, 148535761, 67911621,
              238700391, 224183590, 170998790, 104486975, 81363847, 129161289, 54281363, 100791881,
              185850221, 67400723, 153913781, 247062782, 35411505, 48447796, 90710559, 211284483,
              135389110, 260125445, 26451456, 46126435, 34884345, 199208092, 189299702, 222236846,
              212020732, 157341419, 50385541, 31157387, 214331009, 246555646, 46629005, 38115064,
              200295213, 72618725, 6208689, 145706676, 154135831, 222840723, 99461488, 106939991,
              156023579, 116859647, 47430573, 264758616, 139714595, 184120139, 143466178, 17337072,
              214078274, 38429557, 118216948, 195763450, 264282458, 253615348, 173116375, 3677235,
              197485473, 236609676, 9453674, 126894636, 167134668, 19066791, 157049837, 66528431,
              245518247, 53251080, 43737855, 179997990, 195063937, 41015351, 264289232, 81431484,
              205675156, 64307891, 54092187, 204816575, 251274354, 167135704, 198072981, 91524025,
              44349942, 254723792, 100770703, 75117738, 120419308, 147133292, 224620084, 141917139,
              75240990, 4884476, 267404879, 254692251, 143647295, 124656108, 133881133, 45684920}))
  stage_1_butterfly_1 (
    .x_in(stage_0_per_out[2]),
    .y_in(stage_0_per_out[3]),
    .x_out(stage_1_per_in[2]),
    .y_out(stage_1_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({241419299, 114906207, 189966412, 95956458, 57439678, 93815079, 104968162, 119248786,
              115334054, 244981517, 213018760, 25402945, 66106013, 164849679, 150529015, 253446904,
              66456987, 182759226, 266940341, 65939487, 79732409, 218411001, 61436946, 105651679,
              185097589, 13136617, 230680452, 86425411, 136199054, 248430418, 72619804, 104273059,
              101221270, 48258409, 65241583, 32326785, 161494327, 86611832, 129726580, 248049881,
              227605745, 220409117, 196403691, 60951044, 3059556, 98839404, 262108538, 128923754,
              111262804, 50041017, 39377609, 51590619, 170188367, 71466452, 188624074, 81879124,
              148511346, 6839312, 175901771, 50250252, 109286034, 70993112, 124518160, 202017141,
              40738286, 77785137, 39161232, 166705511, 180106398, 159555178, 219432305, 176106545,
              79909455, 168682489, 259358426, 99151986, 209076586, 45900567, 145040924, 135965343,
              107222748, 95745785, 106026444, 196552678, 136983182, 266184237, 119641299, 36678208,
              231584900, 124689641, 118804291, 250979164, 145952502, 196076822, 58085086, 242448751,
              260055946, 142932928, 26707009, 232700332, 268223107, 26885190, 141552463, 157159811,
              178774268, 187973069, 68124275, 49412866, 5742112, 195777196, 73785583, 24169593,
              186303790, 242906033, 89556414, 123556687, 90238900, 258128862, 211474022, 66398989,
              135620074, 60114085, 80152118, 79759830, 59970273, 203861878, 78067214, 47380903}))
  stage_1_butterfly_2 (
    .x_in(stage_0_per_out[4]),
    .y_in(stage_0_per_out[5]),
    .x_out(stage_1_per_in[4]),
    .y_out(stage_1_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({241419299, 114906207, 189966412, 95956458, 57439678, 93815079, 104968162, 119248786,
              115334054, 244981517, 213018760, 25402945, 66106013, 164849679, 150529015, 253446904,
              66456987, 182759226, 266940341, 65939487, 79732409, 218411001, 61436946, 105651679,
              185097589, 13136617, 230680452, 86425411, 136199054, 248430418, 72619804, 104273059,
              101221270, 48258409, 65241583, 32326785, 161494327, 86611832, 129726580, 248049881,
              227605745, 220409117, 196403691, 60951044, 3059556, 98839404, 262108538, 128923754,
              111262804, 50041017, 39377609, 51590619, 170188367, 71466452, 188624074, 81879124,
              148511346, 6839312, 175901771, 50250252, 109286034, 70993112, 124518160, 202017141,
              40738286, 77785137, 39161232, 166705511, 180106398, 159555178, 219432305, 176106545,
              79909455, 168682489, 259358426, 99151986, 209076586, 45900567, 145040924, 135965343,
              107222748, 95745785, 106026444, 196552678, 136983182, 266184237, 119641299, 36678208,
              231584900, 124689641, 118804291, 250979164, 145952502, 196076822, 58085086, 242448751,
              260055946, 142932928, 26707009, 232700332, 268223107, 26885190, 141552463, 157159811,
              178774268, 187973069, 68124275, 49412866, 5742112, 195777196, 73785583, 24169593,
              186303790, 242906033, 89556414, 123556687, 90238900, 258128862, 211474022, 66398989,
              135620074, 60114085, 80152118, 79759830, 59970273, 203861878, 78067214, 47380903}))
  stage_1_butterfly_3 (
    .x_in(stage_0_per_out[6]),
    .y_in(stage_0_per_out[7]),
    .x_out(stage_1_per_in[6]),
    .y_out(stage_1_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({202037642, 236173805, 141057137, 218922070, 124029413, 59945410, 258951073, 88068083,
              144625416, 184394225, 83042590, 224193580, 152694343, 73580010, 247893310, 38581987,
              113912362, 38792404, 153843002, 22320040, 9977836, 216197112, 203299319, 213462715,
              194834330, 114462613, 127868408, 232970901, 267034870, 264463333, 90431622, 143364478,
              255819997, 127281316, 190155959, 167753662, 92670067, 212643172, 25148713, 182920379,
              10513337, 48499686, 224762304, 145595829, 65501903, 67780496, 72006316, 120068412,
              38583127, 79121294, 138773321, 122372515, 219164507, 4519531, 34739971, 126673466,
              160223263, 233112987, 60791061, 267701123, 202709135, 118263349, 154200425, 83665434,
              111948379, 12994463, 248800534, 106279827, 158020658, 221333762, 20654843, 261080375,
              87171014, 252329804, 84553412, 115935405, 73987125, 205553550, 89839882, 237391515,
              71023991, 154194427, 208367077, 153619107, 109238580, 246502592, 140702439, 248921617,
              144486207, 103784724, 198469359, 96644160, 156384032, 257122505, 243002151, 54591848,
              66619308, 117082039, 255369977, 205764394, 136306850, 85879269, 27101256, 230500375,
              204183192, 91384253, 215044990, 166918201, 37830528, 253166836, 176150397, 58002164,
              230038199, 222792306, 84103703, 174707320, 37832342, 19111856, 109081133, 120623833,
              184194991, 233855133, 161356640, 215876710, 85850918, 74620568, 61148806, 117068649}))
  stage_1_butterfly_4 (
    .x_in(stage_0_per_out[8]),
    .y_in(stage_0_per_out[9]),
    .x_out(stage_1_per_in[8]),
    .y_out(stage_1_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({202037642, 236173805, 141057137, 218922070, 124029413, 59945410, 258951073, 88068083,
              144625416, 184394225, 83042590, 224193580, 152694343, 73580010, 247893310, 38581987,
              113912362, 38792404, 153843002, 22320040, 9977836, 216197112, 203299319, 213462715,
              194834330, 114462613, 127868408, 232970901, 267034870, 264463333, 90431622, 143364478,
              255819997, 127281316, 190155959, 167753662, 92670067, 212643172, 25148713, 182920379,
              10513337, 48499686, 224762304, 145595829, 65501903, 67780496, 72006316, 120068412,
              38583127, 79121294, 138773321, 122372515, 219164507, 4519531, 34739971, 126673466,
              160223263, 233112987, 60791061, 267701123, 202709135, 118263349, 154200425, 83665434,
              111948379, 12994463, 248800534, 106279827, 158020658, 221333762, 20654843, 261080375,
              87171014, 252329804, 84553412, 115935405, 73987125, 205553550, 89839882, 237391515,
              71023991, 154194427, 208367077, 153619107, 109238580, 246502592, 140702439, 248921617,
              144486207, 103784724, 198469359, 96644160, 156384032, 257122505, 243002151, 54591848,
              66619308, 117082039, 255369977, 205764394, 136306850, 85879269, 27101256, 230500375,
              204183192, 91384253, 215044990, 166918201, 37830528, 253166836, 176150397, 58002164,
              230038199, 222792306, 84103703, 174707320, 37832342, 19111856, 109081133, 120623833,
              184194991, 233855133, 161356640, 215876710, 85850918, 74620568, 61148806, 117068649}))
  stage_1_butterfly_5 (
    .x_in(stage_0_per_out[10]),
    .y_in(stage_0_per_out[11]),
    .x_out(stage_1_per_in[10]),
    .y_out(stage_1_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({224076531, 154634100, 75414331, 158913333, 176876579, 195704814, 55709426, 176734838,
              42559975, 100279875, 9179161, 145325214, 181657279, 265093046, 95442771, 11727916,
              179710610, 64402402, 188476710, 60782408, 131815160, 22419281, 214979600, 20002868,
              22106362, 130965208, 127510598, 104683412, 251982020, 239219986, 217412044, 123982174,
              161018204, 185120175, 82911469, 254862428, 54856389, 258398710, 34957318, 86422302,
              141500462, 127264350, 176271587, 95857789, 138344594, 205236983, 207338429, 63759475,
              36505175, 105759020, 35544064, 61255010, 107122996, 65162419, 89363633, 220487343,
              183471966, 199811874, 79351768, 253117467, 263768524, 3615863, 245466834, 114664154,
              79007221, 126437335, 72719897, 78726832, 75051406, 67459976, 104015737, 175735543,
              254205318, 178639438, 77136822, 104494180, 48961458, 43817935, 73243528, 7525756,
              236016875, 219155874, 16967674, 238828812, 41046131, 209365645, 205950205, 21397846,
              263500442, 87333346, 20490089, 59853183, 238066757, 95592544, 176574100, 80415871,
              173525016, 240329350, 215608734, 243959994, 146660836, 83440545, 207179347, 44095704,
              2306944, 109752985, 217413665, 213675734, 233611200, 91771920, 76831465, 83594289,
              249749550, 252048491, 131659808, 215932651, 111544693, 23196483, 252140774, 209775390,
              216035935, 45533578, 201376724, 129973973, 86146205, 153870377, 115561740, 177655074}))
  stage_1_butterfly_6 (
    .x_in(stage_0_per_out[12]),
    .y_in(stage_0_per_out[13]),
    .x_out(stage_1_per_in[12]),
    .y_out(stage_1_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({224076531, 154634100, 75414331, 158913333, 176876579, 195704814, 55709426, 176734838,
              42559975, 100279875, 9179161, 145325214, 181657279, 265093046, 95442771, 11727916,
              179710610, 64402402, 188476710, 60782408, 131815160, 22419281, 214979600, 20002868,
              22106362, 130965208, 127510598, 104683412, 251982020, 239219986, 217412044, 123982174,
              161018204, 185120175, 82911469, 254862428, 54856389, 258398710, 34957318, 86422302,
              141500462, 127264350, 176271587, 95857789, 138344594, 205236983, 207338429, 63759475,
              36505175, 105759020, 35544064, 61255010, 107122996, 65162419, 89363633, 220487343,
              183471966, 199811874, 79351768, 253117467, 263768524, 3615863, 245466834, 114664154,
              79007221, 126437335, 72719897, 78726832, 75051406, 67459976, 104015737, 175735543,
              254205318, 178639438, 77136822, 104494180, 48961458, 43817935, 73243528, 7525756,
              236016875, 219155874, 16967674, 238828812, 41046131, 209365645, 205950205, 21397846,
              263500442, 87333346, 20490089, 59853183, 238066757, 95592544, 176574100, 80415871,
              173525016, 240329350, 215608734, 243959994, 146660836, 83440545, 207179347, 44095704,
              2306944, 109752985, 217413665, 213675734, 233611200, 91771920, 76831465, 83594289,
              249749550, 252048491, 131659808, 215932651, 111544693, 23196483, 252140774, 209775390,
              216035935, 45533578, 201376724, 129973973, 86146205, 153870377, 115561740, 177655074}))
  stage_1_butterfly_7 (
    .x_in(stage_0_per_out[14]),
    .y_in(stage_0_per_out[15]),
    .x_out(stage_1_per_in[14]),
    .y_out(stage_1_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({262853884, 82346526, 204172184, 125480758, 202016934, 58372872, 144194814, 128081279,
              200835165, 226865216, 155441062, 196727396, 139662643, 5284602, 209967729, 133543242,
              213369302, 30998042, 193915015, 53716996, 48721923, 182147827, 222818810, 26713518,
              77445892, 1381761, 151896708, 171508784, 41376169, 57884406, 207289252, 5028136,
              260565899, 126629575, 192679930, 267892175, 80939041, 14425613, 40189829, 50106553,
              28923545, 61366355, 169229772, 14195884, 89821167, 234435452, 74346844, 73917671,
              221852517, 189834774, 216420108, 195995970, 116261862, 193726599, 150921330, 181264550,
              81165688, 224367752, 172134458, 79252444, 254651521, 260962587, 143985240, 125264465,
              251186267, 110001979, 188623776, 264722248, 173013758, 230614882, 192273850, 232215778,
              7373784, 90833651, 202075477, 18807047, 33406019, 41031357, 76213351, 79343207,
              256339290, 223156719, 259641163, 205816155, 2568552, 102404987, 94417879, 192939426,
              66687, 93188095, 82259521, 262718787, 14131216, 95943159, 226423252, 15406607,
              117147237, 216344829, 259932536, 116341913, 2885885, 77043356, 232035425, 148816114,
              69918547, 76840577, 166849602, 145444168, 13809973, 126638229, 217984510, 258312618,
              195258296, 175434645, 144316291, 175360485, 232016200, 228233519, 91036891, 85861280,
              224618046, 21699914, 18026307, 158406994, 24281843, 149817301, 168335279, 146642358}))
  stage_1_butterfly_8 (
    .x_in(stage_0_per_out[16]),
    .y_in(stage_0_per_out[17]),
    .x_out(stage_1_per_in[16]),
    .y_out(stage_1_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({262853884, 82346526, 204172184, 125480758, 202016934, 58372872, 144194814, 128081279,
              200835165, 226865216, 155441062, 196727396, 139662643, 5284602, 209967729, 133543242,
              213369302, 30998042, 193915015, 53716996, 48721923, 182147827, 222818810, 26713518,
              77445892, 1381761, 151896708, 171508784, 41376169, 57884406, 207289252, 5028136,
              260565899, 126629575, 192679930, 267892175, 80939041, 14425613, 40189829, 50106553,
              28923545, 61366355, 169229772, 14195884, 89821167, 234435452, 74346844, 73917671,
              221852517, 189834774, 216420108, 195995970, 116261862, 193726599, 150921330, 181264550,
              81165688, 224367752, 172134458, 79252444, 254651521, 260962587, 143985240, 125264465,
              251186267, 110001979, 188623776, 264722248, 173013758, 230614882, 192273850, 232215778,
              7373784, 90833651, 202075477, 18807047, 33406019, 41031357, 76213351, 79343207,
              256339290, 223156719, 259641163, 205816155, 2568552, 102404987, 94417879, 192939426,
              66687, 93188095, 82259521, 262718787, 14131216, 95943159, 226423252, 15406607,
              117147237, 216344829, 259932536, 116341913, 2885885, 77043356, 232035425, 148816114,
              69918547, 76840577, 166849602, 145444168, 13809973, 126638229, 217984510, 258312618,
              195258296, 175434645, 144316291, 175360485, 232016200, 228233519, 91036891, 85861280,
              224618046, 21699914, 18026307, 158406994, 24281843, 149817301, 168335279, 146642358}))
  stage_1_butterfly_9 (
    .x_in(stage_0_per_out[18]),
    .y_in(stage_0_per_out[19]),
    .x_out(stage_1_per_in[18]),
    .y_out(stage_1_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({243595082, 124972666, 114289273, 59278718, 205274966, 35010964, 80852279, 48487396,
              13214022, 144113751, 183986337, 8772869, 4628244, 146661492, 255259435, 34093582,
              204246510, 248813222, 146691665, 140980229, 27222642, 209335538, 165177241, 264638858,
              90803899, 64059298, 253065021, 187469377, 156486669, 95362545, 182882105, 70333973,
              2705617, 12562435, 171586403, 100306740, 94113816, 121954140, 154399218, 202839194,
              35769351, 133033169, 177621090, 178750844, 180859208, 176649880, 27789608, 132216843,
              234383020, 200991325, 103427147, 203006324, 37907807, 191064173, 180135303, 226857524,
              82858612, 11713205, 111988251, 6515518, 67895486, 24417340, 75455626, 214119665,
              212990958, 50422568, 176645554, 22483780, 239438610, 152117270, 244247525, 52952054,
              82105625, 209487240, 197737960, 119598304, 223749061, 140766862, 204890405, 176646986,
              193207980, 199654780, 258770065, 27342032, 22039584, 237702991, 7487276, 80711179,
              198659369, 53666796, 149046252, 114157546, 33154381, 200880844, 33861678, 184171973,
              46680870, 54194127, 64324001, 104225870, 57534183, 53103748, 212068395, 85943438,
              197375798, 85925921, 248421583, 146917464, 211651639, 39159482, 262436297, 239243318,
              85354678, 82994670, 239135625, 24889364, 230913482, 151554022, 186920055, 165873702,
              242981970, 131606898, 119165597, 71397785, 118812967, 185196127, 88850354, 159375180}))
  stage_1_butterfly_10 (
    .x_in(stage_0_per_out[20]),
    .y_in(stage_0_per_out[21]),
    .x_out(stage_1_per_in[20]),
    .y_out(stage_1_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({243595082, 124972666, 114289273, 59278718, 205274966, 35010964, 80852279, 48487396,
              13214022, 144113751, 183986337, 8772869, 4628244, 146661492, 255259435, 34093582,
              204246510, 248813222, 146691665, 140980229, 27222642, 209335538, 165177241, 264638858,
              90803899, 64059298, 253065021, 187469377, 156486669, 95362545, 182882105, 70333973,
              2705617, 12562435, 171586403, 100306740, 94113816, 121954140, 154399218, 202839194,
              35769351, 133033169, 177621090, 178750844, 180859208, 176649880, 27789608, 132216843,
              234383020, 200991325, 103427147, 203006324, 37907807, 191064173, 180135303, 226857524,
              82858612, 11713205, 111988251, 6515518, 67895486, 24417340, 75455626, 214119665,
              212990958, 50422568, 176645554, 22483780, 239438610, 152117270, 244247525, 52952054,
              82105625, 209487240, 197737960, 119598304, 223749061, 140766862, 204890405, 176646986,
              193207980, 199654780, 258770065, 27342032, 22039584, 237702991, 7487276, 80711179,
              198659369, 53666796, 149046252, 114157546, 33154381, 200880844, 33861678, 184171973,
              46680870, 54194127, 64324001, 104225870, 57534183, 53103748, 212068395, 85943438,
              197375798, 85925921, 248421583, 146917464, 211651639, 39159482, 262436297, 239243318,
              85354678, 82994670, 239135625, 24889364, 230913482, 151554022, 186920055, 165873702,
              242981970, 131606898, 119165597, 71397785, 118812967, 185196127, 88850354, 159375180}))
  stage_1_butterfly_11 (
    .x_in(stage_0_per_out[22]),
    .y_in(stage_0_per_out[23]),
    .x_out(stage_1_per_in[22]),
    .y_out(stage_1_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({256992454, 259902883, 266373219, 64064097, 239354922, 32769539, 34279912, 136417444,
              86047893, 253791818, 209875154, 157208225, 84463383, 90415400, 121172029, 182812696,
              174110644, 141049304, 250769297, 144089543, 116219557, 201671086, 242437879, 81774581,
              35608242, 69255389, 181957723, 256522921, 28513237, 148688834, 25651112, 212200386,
              230880884, 5071752, 207436891, 50115805, 9083394, 18362334, 35697312, 96014882,
              254464819, 134836604, 29380441, 223616593, 63900610, 239800333, 34535827, 241368847,
              37207751, 94872102, 104305160, 38129962, 259466327, 77506253, 22230677, 221869909,
              258848760, 124878920, 245673827, 119697484, 225061179, 163120146, 211697180, 217885801,
              7004663, 96098889, 154780521, 259065776, 156508649, 70871651, 76495986, 41460117,
              193530415, 242696977, 113066699, 25013575, 173627934, 95276657, 112847505, 71010071,
              208392312, 203277373, 139316176, 62424622, 161193348, 28990836, 184571212, 18485653,
              256317058, 16822583, 178875242, 255875272, 96851793, 122635188, 247989601, 155632772,
              104721465, 185121114, 155494097, 134337294, 188253439, 225384963, 147907047, 139206238,
              194631063, 148548934, 243436973, 176530780, 218464636, 41573703, 177240151, 127930513,
              175705236, 231508432, 138028127, 73886338, 144500142, 94729012, 106663692, 52942312,
              250268531, 189935724, 110007683, 75752194, 208182039, 243900215, 78372181, 4980542}))
  stage_1_butterfly_12 (
    .x_in(stage_0_per_out[24]),
    .y_in(stage_0_per_out[25]),
    .x_out(stage_1_per_in[24]),
    .y_out(stage_1_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({256992454, 259902883, 266373219, 64064097, 239354922, 32769539, 34279912, 136417444,
              86047893, 253791818, 209875154, 157208225, 84463383, 90415400, 121172029, 182812696,
              174110644, 141049304, 250769297, 144089543, 116219557, 201671086, 242437879, 81774581,
              35608242, 69255389, 181957723, 256522921, 28513237, 148688834, 25651112, 212200386,
              230880884, 5071752, 207436891, 50115805, 9083394, 18362334, 35697312, 96014882,
              254464819, 134836604, 29380441, 223616593, 63900610, 239800333, 34535827, 241368847,
              37207751, 94872102, 104305160, 38129962, 259466327, 77506253, 22230677, 221869909,
              258848760, 124878920, 245673827, 119697484, 225061179, 163120146, 211697180, 217885801,
              7004663, 96098889, 154780521, 259065776, 156508649, 70871651, 76495986, 41460117,
              193530415, 242696977, 113066699, 25013575, 173627934, 95276657, 112847505, 71010071,
              208392312, 203277373, 139316176, 62424622, 161193348, 28990836, 184571212, 18485653,
              256317058, 16822583, 178875242, 255875272, 96851793, 122635188, 247989601, 155632772,
              104721465, 185121114, 155494097, 134337294, 188253439, 225384963, 147907047, 139206238,
              194631063, 148548934, 243436973, 176530780, 218464636, 41573703, 177240151, 127930513,
              175705236, 231508432, 138028127, 73886338, 144500142, 94729012, 106663692, 52942312,
              250268531, 189935724, 110007683, 75752194, 208182039, 243900215, 78372181, 4980542}))
  stage_1_butterfly_13 (
    .x_in(stage_0_per_out[26]),
    .y_in(stage_0_per_out[27]),
    .x_out(stage_1_per_in[26]),
    .y_out(stage_1_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({77239454, 127717239, 148884778, 135644103, 143734200, 6456449, 236741674, 157158700,
              222855093, 172630653, 57044952, 51299486, 86334506, 217483488, 126959268, 254780782,
              21923530, 137520333, 126650083, 50213981, 186026798, 139730465, 33343400, 108532653,
              26776855, 248206642, 40931981, 34242638, 42903438, 22116392, 63912782, 134518349,
              58103200, 259334239, 166350047, 152505970, 239780428, 13394971, 91136142, 187892585,
              251689720, 112174110, 110850189, 254241553, 253128696, 179888950, 81924749, 256890018,
              197145719, 16703359, 187446019, 35688570, 56848151, 197641184, 255364493, 153805373,
              164222678, 143389876, 124441328, 258225039, 79432680, 74661667, 39292866, 50021352,
              143288167, 75588758, 210949816, 209423491, 22021280, 4184358, 117619035, 179675005,
              248341796, 33161823, 123481104, 31515852, 27523605, 107466416, 153827860, 244217621,
              197016099, 14369566, 250734390, 27456585, 171258656, 243789725, 106713399, 94477870,
              262755833, 133797547, 108936038, 207692352, 60493834, 38723858, 152193297, 12048336,
              13327732, 227177249, 130184658, 48893661, 14594411, 215351473, 260941520, 102888853,
              193102647, 55952036, 267667077, 157311612, 218565763, 192111834, 162889363, 116226,
              57880935, 186728485, 98151275, 187345691, 202657965, 153057061, 141192231, 106441080,
              145663803, 170437415, 142379740, 126420356, 68372869, 6554463, 252921174, 101380813}))
  stage_1_butterfly_14 (
    .x_in(stage_0_per_out[28]),
    .y_in(stage_0_per_out[29]),
    .x_out(stage_1_per_in[28]),
    .y_out(stage_1_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[1]),
    .factors({77239454, 127717239, 148884778, 135644103, 143734200, 6456449, 236741674, 157158700,
              222855093, 172630653, 57044952, 51299486, 86334506, 217483488, 126959268, 254780782,
              21923530, 137520333, 126650083, 50213981, 186026798, 139730465, 33343400, 108532653,
              26776855, 248206642, 40931981, 34242638, 42903438, 22116392, 63912782, 134518349,
              58103200, 259334239, 166350047, 152505970, 239780428, 13394971, 91136142, 187892585,
              251689720, 112174110, 110850189, 254241553, 253128696, 179888950, 81924749, 256890018,
              197145719, 16703359, 187446019, 35688570, 56848151, 197641184, 255364493, 153805373,
              164222678, 143389876, 124441328, 258225039, 79432680, 74661667, 39292866, 50021352,
              143288167, 75588758, 210949816, 209423491, 22021280, 4184358, 117619035, 179675005,
              248341796, 33161823, 123481104, 31515852, 27523605, 107466416, 153827860, 244217621,
              197016099, 14369566, 250734390, 27456585, 171258656, 243789725, 106713399, 94477870,
              262755833, 133797547, 108936038, 207692352, 60493834, 38723858, 152193297, 12048336,
              13327732, 227177249, 130184658, 48893661, 14594411, 215351473, 260941520, 102888853,
              193102647, 55952036, 267667077, 157311612, 218565763, 192111834, 162889363, 116226,
              57880935, 186728485, 98151275, 187345691, 202657965, 153057061, 141192231, 106441080,
              145663803, 170437415, 142379740, 126420356, 68372869, 6554463, 252921174, 101380813}))
  stage_1_butterfly_15 (
    .x_in(stage_0_per_out[30]),
    .y_in(stage_0_per_out[31]),
    .x_out(stage_1_per_in[30]),
    .y_out(stage_1_per_in[31]),
    .clk(clk),
    .rst(rst)
  );




  
  // TODO(Yang): stage 1 -> stage 2 permutation
  // FIXME: ignore butterfly units for now.
  stage_1_permutation #(
    .DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    .INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_1_2_per (
    .inData_0(stage_1_per_in[0]),
    .inData_1(stage_1_per_in[1]),
    .inData_2(stage_1_per_in[2]),
    .inData_3(stage_1_per_in[3]),
    .inData_4(stage_1_per_in[4]),
    .inData_5(stage_1_per_in[5]),
    .inData_6(stage_1_per_in[6]),
    .inData_7(stage_1_per_in[7]),
    .inData_8(stage_1_per_in[8]),
    .inData_9(stage_1_per_in[9]),
    .inData_10(stage_1_per_in[10]),
    .inData_11(stage_1_per_in[11]),
    .inData_12(stage_1_per_in[12]),
    .inData_13(stage_1_per_in[13]),
    .inData_14(stage_1_per_in[14]),
    .inData_15(stage_1_per_in[15]),
    .inData_16(stage_1_per_in[16]),
    .inData_17(stage_1_per_in[17]),
    .inData_18(stage_1_per_in[18]),
    .inData_19(stage_1_per_in[19]),
    .inData_20(stage_1_per_in[20]),
    .inData_21(stage_1_per_in[21]),
    .inData_22(stage_1_per_in[22]),
    .inData_23(stage_1_per_in[23]),
    .inData_24(stage_1_per_in[24]),
    .inData_25(stage_1_per_in[25]),
    .inData_26(stage_1_per_in[26]),
    .inData_27(stage_1_per_in[27]),
    .inData_28(stage_1_per_in[28]),
    .inData_29(stage_1_per_in[29]),
    .inData_30(stage_1_per_in[30]),
    .inData_31(stage_1_per_in[31]),
    .outData_0(stage_1_per_out[0]),
    .outData_1(stage_1_per_out[1]),
    .outData_2(stage_1_per_out[2]),
    .outData_3(stage_1_per_out[3]),
    .outData_4(stage_1_per_out[4]),
    .outData_5(stage_1_per_out[5]),
    .outData_6(stage_1_per_out[6]),
    .outData_7(stage_1_per_out[7]),
    .outData_8(stage_1_per_out[8]),
    .outData_9(stage_1_per_out[9]),
    .outData_10(stage_1_per_out[10]),
    .outData_11(stage_1_per_out[11]),
    .outData_12(stage_1_per_out[12]),
    .outData_13(stage_1_per_out[13]),
    .outData_14(stage_1_per_out[14]),
    .outData_15(stage_1_per_out[15]),
    .outData_16(stage_1_per_out[16]),
    .outData_17(stage_1_per_out[17]),
    .outData_18(stage_1_per_out[18]),
    .outData_19(stage_1_per_out[19]),
    .outData_20(stage_1_per_out[20]),
    .outData_21(stage_1_per_out[21]),
    .outData_22(stage_1_per_out[22]),
    .outData_23(stage_1_per_out[23]),
    .outData_24(stage_1_per_out[24]),
    .outData_25(stage_1_per_out[25]),
    .outData_26(stage_1_per_out[26]),
    .outData_27(stage_1_per_out[27]),
    .outData_28(stage_1_per_out[28]),
    .outData_29(stage_1_per_out[29]),
    .outData_30(stage_1_per_out[30]),
    .outData_31(stage_1_per_out[31]),
    .in_start(in_start[1]),
    .out_start(out_start[1]),
    .clk(clk),
    .rst(rst)
  );


  // TODO(Tian): stage 2 32 butterfly units
  butterfly #(
    .start(START_CYCLE[2]),
    .factors({187381670, 64830196, 235273242, 266562472, 120217110, 70325928, 135902522, 232847226,
              54714468, 163197321, 249576229, 83977288, 142656304, 102034957, 122969043, 144502563,
              196018390, 31964447, 206341936, 262112169, 212112171, 251717800, 81414740, 107503597,
              26068775, 9205704, 141956852, 217359458, 174191574, 85566308, 209112367, 184177651,
              27439037, 148108490, 72369588, 172401093, 189139684, 237616434, 265348407, 5161923,
              58661398, 128052734, 1855205, 22997488, 128297265, 113049121, 171206517, 252018541,
              174612628, 261143222, 226834391, 584543, 23442787, 211201491, 77127228, 183571221,
              35629855, 151857114, 43000087, 198336839, 50083600, 53025186, 246787643, 66582189,
              233083676, 74918627, 237125965, 142807968, 24365404, 83194655, 244423105, 174290656,
              173628384, 31540722, 85740049, 87492030, 63661975, 167181901, 90687088, 22383105,
              142941966, 32160642, 167645260, 46312994, 252714435, 38415865, 145831337, 238775640,
              10646661, 264974639, 206116619, 248328138, 156195364, 36213609, 191744986, 250611881,
              250031819, 156534179, 121730405, 209698557, 183613005, 148649408, 205856513, 227453822,
              206844979, 42575603, 174028560, 93513491, 78273516, 263102666, 175598948, 169092523,
              121414397, 47531240, 4721397, 258059551, 72509307, 212425161, 146344523, 139742686,
              255478273, 19817676, 62435894, 131659168, 255463943, 25652741, 193174373, 113269084}))
  stage_2_butterfly_0 (
    .x_in(stage_1_per_out[0]),
    .y_in(stage_1_per_out[1]),
    .x_out(stage_2_per_in[0]),
    .y_out(stage_2_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({187381670, 64830196, 235273242, 266562472, 120217110, 70325928, 135902522, 232847226,
              54714468, 163197321, 249576229, 83977288, 142656304, 102034957, 122969043, 144502563,
              196018390, 31964447, 206341936, 262112169, 212112171, 251717800, 81414740, 107503597,
              26068775, 9205704, 141956852, 217359458, 174191574, 85566308, 209112367, 184177651,
              27439037, 148108490, 72369588, 172401093, 189139684, 237616434, 265348407, 5161923,
              58661398, 128052734, 1855205, 22997488, 128297265, 113049121, 171206517, 252018541,
              174612628, 261143222, 226834391, 584543, 23442787, 211201491, 77127228, 183571221,
              35629855, 151857114, 43000087, 198336839, 50083600, 53025186, 246787643, 66582189,
              233083676, 74918627, 237125965, 142807968, 24365404, 83194655, 244423105, 174290656,
              173628384, 31540722, 85740049, 87492030, 63661975, 167181901, 90687088, 22383105,
              142941966, 32160642, 167645260, 46312994, 252714435, 38415865, 145831337, 238775640,
              10646661, 264974639, 206116619, 248328138, 156195364, 36213609, 191744986, 250611881,
              250031819, 156534179, 121730405, 209698557, 183613005, 148649408, 205856513, 227453822,
              206844979, 42575603, 174028560, 93513491, 78273516, 263102666, 175598948, 169092523,
              121414397, 47531240, 4721397, 258059551, 72509307, 212425161, 146344523, 139742686,
              255478273, 19817676, 62435894, 131659168, 255463943, 25652741, 193174373, 113269084}))
  stage_2_butterfly_1 (
    .x_in(stage_1_per_out[2]),
    .y_in(stage_1_per_out[3]),
    .x_out(stage_2_per_in[2]),
    .y_out(stage_2_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({187381670, 64830196, 235273242, 266562472, 120217110, 70325928, 135902522, 232847226,
              54714468, 163197321, 249576229, 83977288, 142656304, 102034957, 122969043, 144502563,
              196018390, 31964447, 206341936, 262112169, 212112171, 251717800, 81414740, 107503597,
              26068775, 9205704, 141956852, 217359458, 174191574, 85566308, 209112367, 184177651,
              27439037, 148108490, 72369588, 172401093, 189139684, 237616434, 265348407, 5161923,
              58661398, 128052734, 1855205, 22997488, 128297265, 113049121, 171206517, 252018541,
              174612628, 261143222, 226834391, 584543, 23442787, 211201491, 77127228, 183571221,
              35629855, 151857114, 43000087, 198336839, 50083600, 53025186, 246787643, 66582189,
              233083676, 74918627, 237125965, 142807968, 24365404, 83194655, 244423105, 174290656,
              173628384, 31540722, 85740049, 87492030, 63661975, 167181901, 90687088, 22383105,
              142941966, 32160642, 167645260, 46312994, 252714435, 38415865, 145831337, 238775640,
              10646661, 264974639, 206116619, 248328138, 156195364, 36213609, 191744986, 250611881,
              250031819, 156534179, 121730405, 209698557, 183613005, 148649408, 205856513, 227453822,
              206844979, 42575603, 174028560, 93513491, 78273516, 263102666, 175598948, 169092523,
              121414397, 47531240, 4721397, 258059551, 72509307, 212425161, 146344523, 139742686,
              255478273, 19817676, 62435894, 131659168, 255463943, 25652741, 193174373, 113269084}))
  stage_2_butterfly_2 (
    .x_in(stage_1_per_out[4]),
    .y_in(stage_1_per_out[5]),
    .x_out(stage_2_per_in[4]),
    .y_out(stage_2_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({187381670, 64830196, 235273242, 266562472, 120217110, 70325928, 135902522, 232847226,
              54714468, 163197321, 249576229, 83977288, 142656304, 102034957, 122969043, 144502563,
              196018390, 31964447, 206341936, 262112169, 212112171, 251717800, 81414740, 107503597,
              26068775, 9205704, 141956852, 217359458, 174191574, 85566308, 209112367, 184177651,
              27439037, 148108490, 72369588, 172401093, 189139684, 237616434, 265348407, 5161923,
              58661398, 128052734, 1855205, 22997488, 128297265, 113049121, 171206517, 252018541,
              174612628, 261143222, 226834391, 584543, 23442787, 211201491, 77127228, 183571221,
              35629855, 151857114, 43000087, 198336839, 50083600, 53025186, 246787643, 66582189,
              233083676, 74918627, 237125965, 142807968, 24365404, 83194655, 244423105, 174290656,
              173628384, 31540722, 85740049, 87492030, 63661975, 167181901, 90687088, 22383105,
              142941966, 32160642, 167645260, 46312994, 252714435, 38415865, 145831337, 238775640,
              10646661, 264974639, 206116619, 248328138, 156195364, 36213609, 191744986, 250611881,
              250031819, 156534179, 121730405, 209698557, 183613005, 148649408, 205856513, 227453822,
              206844979, 42575603, 174028560, 93513491, 78273516, 263102666, 175598948, 169092523,
              121414397, 47531240, 4721397, 258059551, 72509307, 212425161, 146344523, 139742686,
              255478273, 19817676, 62435894, 131659168, 255463943, 25652741, 193174373, 113269084}))
  stage_2_butterfly_3 (
    .x_in(stage_1_per_out[6]),
    .y_in(stage_1_per_out[7]),
    .x_out(stage_2_per_in[6]),
    .y_out(stage_2_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({222912429, 62456195, 77536776, 65498827, 248922055, 139101859, 189601976, 181593250,
              38252193, 18205961, 155363318, 73685379, 157839041, 107513427, 94792077, 133098101,
              243009216, 90701762, 65889055, 245041907, 21649526, 228715598, 164248031, 133952844,
              187208958, 122609533, 212237706, 69412414, 116527240, 37504237, 261541195, 149904904,
              189909138, 157649589, 205242220, 265496406, 190586128, 102785717, 34052825, 55947412,
              224322272, 123720956, 86359417, 134561032, 130154791, 212728405, 254842567, 131471427,
              75993973, 163812077, 169792793, 228572460, 259621463, 257402730, 146205579, 121970089,
              509728, 29537138, 256834872, 186476418, 190565686, 248946430, 159538295, 120318911,
              82779345, 129694458, 250727821, 149925004, 211982342, 222087036, 243339369, 236528116,
              58491201, 183590673, 56723699, 210373784, 147903734, 111532362, 224922683, 53126225,
              128589211, 12711531, 191250025, 137060289, 165001005, 162575967, 136179523, 255737752,
              267008435, 86752434, 61322741, 4457103, 147014646, 153316076, 57946842, 157386503,
              54690936, 61348732, 100611174, 23776027, 174163034, 67784869, 56545684, 212162524,
              53284215, 168674209, 148479452, 203905228, 226025718, 199055975, 161217010, 50376784,
              156298941, 5368199, 141267184, 203598031, 73072346, 37377133, 5739737, 134804553,
              186048173, 127918992, 223481427, 193897399, 112360014, 143811089, 103896237, 149423455}))
  stage_2_butterfly_4 (
    .x_in(stage_1_per_out[8]),
    .y_in(stage_1_per_out[9]),
    .x_out(stage_2_per_in[8]),
    .y_out(stage_2_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({222912429, 62456195, 77536776, 65498827, 248922055, 139101859, 189601976, 181593250,
              38252193, 18205961, 155363318, 73685379, 157839041, 107513427, 94792077, 133098101,
              243009216, 90701762, 65889055, 245041907, 21649526, 228715598, 164248031, 133952844,
              187208958, 122609533, 212237706, 69412414, 116527240, 37504237, 261541195, 149904904,
              189909138, 157649589, 205242220, 265496406, 190586128, 102785717, 34052825, 55947412,
              224322272, 123720956, 86359417, 134561032, 130154791, 212728405, 254842567, 131471427,
              75993973, 163812077, 169792793, 228572460, 259621463, 257402730, 146205579, 121970089,
              509728, 29537138, 256834872, 186476418, 190565686, 248946430, 159538295, 120318911,
              82779345, 129694458, 250727821, 149925004, 211982342, 222087036, 243339369, 236528116,
              58491201, 183590673, 56723699, 210373784, 147903734, 111532362, 224922683, 53126225,
              128589211, 12711531, 191250025, 137060289, 165001005, 162575967, 136179523, 255737752,
              267008435, 86752434, 61322741, 4457103, 147014646, 153316076, 57946842, 157386503,
              54690936, 61348732, 100611174, 23776027, 174163034, 67784869, 56545684, 212162524,
              53284215, 168674209, 148479452, 203905228, 226025718, 199055975, 161217010, 50376784,
              156298941, 5368199, 141267184, 203598031, 73072346, 37377133, 5739737, 134804553,
              186048173, 127918992, 223481427, 193897399, 112360014, 143811089, 103896237, 149423455}))
  stage_2_butterfly_5 (
    .x_in(stage_1_per_out[10]),
    .y_in(stage_1_per_out[11]),
    .x_out(stage_2_per_in[10]),
    .y_out(stage_2_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({222912429, 62456195, 77536776, 65498827, 248922055, 139101859, 189601976, 181593250,
              38252193, 18205961, 155363318, 73685379, 157839041, 107513427, 94792077, 133098101,
              243009216, 90701762, 65889055, 245041907, 21649526, 228715598, 164248031, 133952844,
              187208958, 122609533, 212237706, 69412414, 116527240, 37504237, 261541195, 149904904,
              189909138, 157649589, 205242220, 265496406, 190586128, 102785717, 34052825, 55947412,
              224322272, 123720956, 86359417, 134561032, 130154791, 212728405, 254842567, 131471427,
              75993973, 163812077, 169792793, 228572460, 259621463, 257402730, 146205579, 121970089,
              509728, 29537138, 256834872, 186476418, 190565686, 248946430, 159538295, 120318911,
              82779345, 129694458, 250727821, 149925004, 211982342, 222087036, 243339369, 236528116,
              58491201, 183590673, 56723699, 210373784, 147903734, 111532362, 224922683, 53126225,
              128589211, 12711531, 191250025, 137060289, 165001005, 162575967, 136179523, 255737752,
              267008435, 86752434, 61322741, 4457103, 147014646, 153316076, 57946842, 157386503,
              54690936, 61348732, 100611174, 23776027, 174163034, 67784869, 56545684, 212162524,
              53284215, 168674209, 148479452, 203905228, 226025718, 199055975, 161217010, 50376784,
              156298941, 5368199, 141267184, 203598031, 73072346, 37377133, 5739737, 134804553,
              186048173, 127918992, 223481427, 193897399, 112360014, 143811089, 103896237, 149423455}))
  stage_2_butterfly_6 (
    .x_in(stage_1_per_out[12]),
    .y_in(stage_1_per_out[13]),
    .x_out(stage_2_per_in[12]),
    .y_out(stage_2_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({222912429, 62456195, 77536776, 65498827, 248922055, 139101859, 189601976, 181593250,
              38252193, 18205961, 155363318, 73685379, 157839041, 107513427, 94792077, 133098101,
              243009216, 90701762, 65889055, 245041907, 21649526, 228715598, 164248031, 133952844,
              187208958, 122609533, 212237706, 69412414, 116527240, 37504237, 261541195, 149904904,
              189909138, 157649589, 205242220, 265496406, 190586128, 102785717, 34052825, 55947412,
              224322272, 123720956, 86359417, 134561032, 130154791, 212728405, 254842567, 131471427,
              75993973, 163812077, 169792793, 228572460, 259621463, 257402730, 146205579, 121970089,
              509728, 29537138, 256834872, 186476418, 190565686, 248946430, 159538295, 120318911,
              82779345, 129694458, 250727821, 149925004, 211982342, 222087036, 243339369, 236528116,
              58491201, 183590673, 56723699, 210373784, 147903734, 111532362, 224922683, 53126225,
              128589211, 12711531, 191250025, 137060289, 165001005, 162575967, 136179523, 255737752,
              267008435, 86752434, 61322741, 4457103, 147014646, 153316076, 57946842, 157386503,
              54690936, 61348732, 100611174, 23776027, 174163034, 67784869, 56545684, 212162524,
              53284215, 168674209, 148479452, 203905228, 226025718, 199055975, 161217010, 50376784,
              156298941, 5368199, 141267184, 203598031, 73072346, 37377133, 5739737, 134804553,
              186048173, 127918992, 223481427, 193897399, 112360014, 143811089, 103896237, 149423455}))
  stage_2_butterfly_7 (
    .x_in(stage_1_per_out[14]),
    .y_in(stage_1_per_out[15]),
    .x_out(stage_2_per_in[14]),
    .y_out(stage_2_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({224391994, 48885659, 73481957, 98410858, 29779638, 205681680, 116513948, 16697663,
              217763430, 46120362, 89028484, 163823140, 107830842, 175949223, 187106042, 56081948,
              193911793, 233437339, 207877484, 121712648, 168470500, 127163336, 58903295, 53432143,
              267506256, 79843127, 12286825, 265883664, 82483914, 90149574, 77916555, 94856770,
              231354349, 158914825, 181167176, 126807666, 133273987, 248133554, 145351880, 23586243,
              149788353, 264322432, 160204962, 123313741, 6760936, 229032903, 45355620, 232038388,
              54916848, 7376627, 129325164, 217846048, 207530748, 4643973, 259302720, 106743034,
              36492987, 120080647, 51550886, 121145061, 91458750, 98269185, 110378476, 2487567,
              202032572, 92379159, 218380292, 6001670, 69017626, 160048836, 140358303, 55581691,
              139374293, 184522009, 3260661, 170230234, 268043824, 254234203, 19058782, 180764097,
              158314046, 100343421, 190540901, 103503994, 121608761, 195181845, 222527593, 37498403,
              153237233, 66412546, 60600589, 99996719, 159491687, 126749676, 202565947, 5445105,
              19700796, 247452694, 50174239, 62094530, 8474832, 266777211, 226759664, 219133933,
              81838336, 12551837, 46197346, 55222727, 148491526, 161345834, 92902456, 183669067,
              13228372, 255457916, 78552959, 263649093, 255552842, 59214954, 159148996, 101579460,
              8836114, 110302060, 76313029, 7301415, 256519333, 135080569, 24036023, 168342750}))
  stage_2_butterfly_8 (
    .x_in(stage_1_per_out[16]),
    .y_in(stage_1_per_out[17]),
    .x_out(stage_2_per_in[16]),
    .y_out(stage_2_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({224391994, 48885659, 73481957, 98410858, 29779638, 205681680, 116513948, 16697663,
              217763430, 46120362, 89028484, 163823140, 107830842, 175949223, 187106042, 56081948,
              193911793, 233437339, 207877484, 121712648, 168470500, 127163336, 58903295, 53432143,
              267506256, 79843127, 12286825, 265883664, 82483914, 90149574, 77916555, 94856770,
              231354349, 158914825, 181167176, 126807666, 133273987, 248133554, 145351880, 23586243,
              149788353, 264322432, 160204962, 123313741, 6760936, 229032903, 45355620, 232038388,
              54916848, 7376627, 129325164, 217846048, 207530748, 4643973, 259302720, 106743034,
              36492987, 120080647, 51550886, 121145061, 91458750, 98269185, 110378476, 2487567,
              202032572, 92379159, 218380292, 6001670, 69017626, 160048836, 140358303, 55581691,
              139374293, 184522009, 3260661, 170230234, 268043824, 254234203, 19058782, 180764097,
              158314046, 100343421, 190540901, 103503994, 121608761, 195181845, 222527593, 37498403,
              153237233, 66412546, 60600589, 99996719, 159491687, 126749676, 202565947, 5445105,
              19700796, 247452694, 50174239, 62094530, 8474832, 266777211, 226759664, 219133933,
              81838336, 12551837, 46197346, 55222727, 148491526, 161345834, 92902456, 183669067,
              13228372, 255457916, 78552959, 263649093, 255552842, 59214954, 159148996, 101579460,
              8836114, 110302060, 76313029, 7301415, 256519333, 135080569, 24036023, 168342750}))
  stage_2_butterfly_9 (
    .x_in(stage_1_per_out[18]),
    .y_in(stage_1_per_out[19]),
    .x_out(stage_2_per_in[18]),
    .y_out(stage_2_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({224391994, 48885659, 73481957, 98410858, 29779638, 205681680, 116513948, 16697663,
              217763430, 46120362, 89028484, 163823140, 107830842, 175949223, 187106042, 56081948,
              193911793, 233437339, 207877484, 121712648, 168470500, 127163336, 58903295, 53432143,
              267506256, 79843127, 12286825, 265883664, 82483914, 90149574, 77916555, 94856770,
              231354349, 158914825, 181167176, 126807666, 133273987, 248133554, 145351880, 23586243,
              149788353, 264322432, 160204962, 123313741, 6760936, 229032903, 45355620, 232038388,
              54916848, 7376627, 129325164, 217846048, 207530748, 4643973, 259302720, 106743034,
              36492987, 120080647, 51550886, 121145061, 91458750, 98269185, 110378476, 2487567,
              202032572, 92379159, 218380292, 6001670, 69017626, 160048836, 140358303, 55581691,
              139374293, 184522009, 3260661, 170230234, 268043824, 254234203, 19058782, 180764097,
              158314046, 100343421, 190540901, 103503994, 121608761, 195181845, 222527593, 37498403,
              153237233, 66412546, 60600589, 99996719, 159491687, 126749676, 202565947, 5445105,
              19700796, 247452694, 50174239, 62094530, 8474832, 266777211, 226759664, 219133933,
              81838336, 12551837, 46197346, 55222727, 148491526, 161345834, 92902456, 183669067,
              13228372, 255457916, 78552959, 263649093, 255552842, 59214954, 159148996, 101579460,
              8836114, 110302060, 76313029, 7301415, 256519333, 135080569, 24036023, 168342750}))
  stage_2_butterfly_10 (
    .x_in(stage_1_per_out[20]),
    .y_in(stage_1_per_out[21]),
    .x_out(stage_2_per_in[20]),
    .y_out(stage_2_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({224391994, 48885659, 73481957, 98410858, 29779638, 205681680, 116513948, 16697663,
              217763430, 46120362, 89028484, 163823140, 107830842, 175949223, 187106042, 56081948,
              193911793, 233437339, 207877484, 121712648, 168470500, 127163336, 58903295, 53432143,
              267506256, 79843127, 12286825, 265883664, 82483914, 90149574, 77916555, 94856770,
              231354349, 158914825, 181167176, 126807666, 133273987, 248133554, 145351880, 23586243,
              149788353, 264322432, 160204962, 123313741, 6760936, 229032903, 45355620, 232038388,
              54916848, 7376627, 129325164, 217846048, 207530748, 4643973, 259302720, 106743034,
              36492987, 120080647, 51550886, 121145061, 91458750, 98269185, 110378476, 2487567,
              202032572, 92379159, 218380292, 6001670, 69017626, 160048836, 140358303, 55581691,
              139374293, 184522009, 3260661, 170230234, 268043824, 254234203, 19058782, 180764097,
              158314046, 100343421, 190540901, 103503994, 121608761, 195181845, 222527593, 37498403,
              153237233, 66412546, 60600589, 99996719, 159491687, 126749676, 202565947, 5445105,
              19700796, 247452694, 50174239, 62094530, 8474832, 266777211, 226759664, 219133933,
              81838336, 12551837, 46197346, 55222727, 148491526, 161345834, 92902456, 183669067,
              13228372, 255457916, 78552959, 263649093, 255552842, 59214954, 159148996, 101579460,
              8836114, 110302060, 76313029, 7301415, 256519333, 135080569, 24036023, 168342750}))
  stage_2_butterfly_11 (
    .x_in(stage_1_per_out[22]),
    .y_in(stage_1_per_out[23]),
    .x_out(stage_2_per_in[22]),
    .y_out(stage_2_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({134161265, 2017030, 183700349, 217210388, 165671105, 166139329, 188535281, 17682401,
              184464011, 20118393, 174391063, 60051251, 218207344, 112756762, 266378632, 107138937,
              236272786, 95713937, 150049787, 209744644, 33594840, 224550271, 189044804, 86350556,
              197065781, 67209795, 175710456, 112825183, 14882191, 248465751, 104215821, 24347842,
              114052864, 216531417, 159987098, 62765404, 129677075, 171841734, 140210175, 19637177,
              189757297, 10943590, 72677507, 81197166, 159978713, 7280660, 197425604, 244216061,
              171198428, 267017218, 92441360, 223473865, 195152646, 105443909, 58726750, 29901564,
              99543252, 154298223, 236050384, 160429892, 94436408, 247116469, 153319834, 30998914,
              36196902, 227628318, 135921552, 102243739, 160050812, 138513718, 161607031, 21628090,
              20655050, 166586238, 9793208, 226981541, 145034434, 75689102, 52844710, 95654178,
              233967292, 195298807, 69205492, 198352904, 134796549, 266777383, 187867192, 189248215,
              184560259, 265028258, 164728317, 103189081, 99012968, 151297332, 243091016, 231749609,
              243047656, 228243008, 8650362, 58589536, 54393228, 104290760, 8259535, 74931497,
              94686133, 67241659, 79336225, 255778637, 195270185, 176972907, 234786570, 178382895,
              249947221, 116257755, 123052007, 80381167, 132747224, 27298769, 261458154, 203850982,
              237395333, 122455193, 129740611, 18433789, 227454343, 208475153, 2204580, 98445813}))
  stage_2_butterfly_12 (
    .x_in(stage_1_per_out[24]),
    .y_in(stage_1_per_out[25]),
    .x_out(stage_2_per_in[24]),
    .y_out(stage_2_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({134161265, 2017030, 183700349, 217210388, 165671105, 166139329, 188535281, 17682401,
              184464011, 20118393, 174391063, 60051251, 218207344, 112756762, 266378632, 107138937,
              236272786, 95713937, 150049787, 209744644, 33594840, 224550271, 189044804, 86350556,
              197065781, 67209795, 175710456, 112825183, 14882191, 248465751, 104215821, 24347842,
              114052864, 216531417, 159987098, 62765404, 129677075, 171841734, 140210175, 19637177,
              189757297, 10943590, 72677507, 81197166, 159978713, 7280660, 197425604, 244216061,
              171198428, 267017218, 92441360, 223473865, 195152646, 105443909, 58726750, 29901564,
              99543252, 154298223, 236050384, 160429892, 94436408, 247116469, 153319834, 30998914,
              36196902, 227628318, 135921552, 102243739, 160050812, 138513718, 161607031, 21628090,
              20655050, 166586238, 9793208, 226981541, 145034434, 75689102, 52844710, 95654178,
              233967292, 195298807, 69205492, 198352904, 134796549, 266777383, 187867192, 189248215,
              184560259, 265028258, 164728317, 103189081, 99012968, 151297332, 243091016, 231749609,
              243047656, 228243008, 8650362, 58589536, 54393228, 104290760, 8259535, 74931497,
              94686133, 67241659, 79336225, 255778637, 195270185, 176972907, 234786570, 178382895,
              249947221, 116257755, 123052007, 80381167, 132747224, 27298769, 261458154, 203850982,
              237395333, 122455193, 129740611, 18433789, 227454343, 208475153, 2204580, 98445813}))
  stage_2_butterfly_13 (
    .x_in(stage_1_per_out[26]),
    .y_in(stage_1_per_out[27]),
    .x_out(stage_2_per_in[26]),
    .y_out(stage_2_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({134161265, 2017030, 183700349, 217210388, 165671105, 166139329, 188535281, 17682401,
              184464011, 20118393, 174391063, 60051251, 218207344, 112756762, 266378632, 107138937,
              236272786, 95713937, 150049787, 209744644, 33594840, 224550271, 189044804, 86350556,
              197065781, 67209795, 175710456, 112825183, 14882191, 248465751, 104215821, 24347842,
              114052864, 216531417, 159987098, 62765404, 129677075, 171841734, 140210175, 19637177,
              189757297, 10943590, 72677507, 81197166, 159978713, 7280660, 197425604, 244216061,
              171198428, 267017218, 92441360, 223473865, 195152646, 105443909, 58726750, 29901564,
              99543252, 154298223, 236050384, 160429892, 94436408, 247116469, 153319834, 30998914,
              36196902, 227628318, 135921552, 102243739, 160050812, 138513718, 161607031, 21628090,
              20655050, 166586238, 9793208, 226981541, 145034434, 75689102, 52844710, 95654178,
              233967292, 195298807, 69205492, 198352904, 134796549, 266777383, 187867192, 189248215,
              184560259, 265028258, 164728317, 103189081, 99012968, 151297332, 243091016, 231749609,
              243047656, 228243008, 8650362, 58589536, 54393228, 104290760, 8259535, 74931497,
              94686133, 67241659, 79336225, 255778637, 195270185, 176972907, 234786570, 178382895,
              249947221, 116257755, 123052007, 80381167, 132747224, 27298769, 261458154, 203850982,
              237395333, 122455193, 129740611, 18433789, 227454343, 208475153, 2204580, 98445813}))
  stage_2_butterfly_14 (
    .x_in(stage_1_per_out[28]),
    .y_in(stage_1_per_out[29]),
    .x_out(stage_2_per_in[28]),
    .y_out(stage_2_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[2]),
    .factors({134161265, 2017030, 183700349, 217210388, 165671105, 166139329, 188535281, 17682401,
              184464011, 20118393, 174391063, 60051251, 218207344, 112756762, 266378632, 107138937,
              236272786, 95713937, 150049787, 209744644, 33594840, 224550271, 189044804, 86350556,
              197065781, 67209795, 175710456, 112825183, 14882191, 248465751, 104215821, 24347842,
              114052864, 216531417, 159987098, 62765404, 129677075, 171841734, 140210175, 19637177,
              189757297, 10943590, 72677507, 81197166, 159978713, 7280660, 197425604, 244216061,
              171198428, 267017218, 92441360, 223473865, 195152646, 105443909, 58726750, 29901564,
              99543252, 154298223, 236050384, 160429892, 94436408, 247116469, 153319834, 30998914,
              36196902, 227628318, 135921552, 102243739, 160050812, 138513718, 161607031, 21628090,
              20655050, 166586238, 9793208, 226981541, 145034434, 75689102, 52844710, 95654178,
              233967292, 195298807, 69205492, 198352904, 134796549, 266777383, 187867192, 189248215,
              184560259, 265028258, 164728317, 103189081, 99012968, 151297332, 243091016, 231749609,
              243047656, 228243008, 8650362, 58589536, 54393228, 104290760, 8259535, 74931497,
              94686133, 67241659, 79336225, 255778637, 195270185, 176972907, 234786570, 178382895,
              249947221, 116257755, 123052007, 80381167, 132747224, 27298769, 261458154, 203850982,
              237395333, 122455193, 129740611, 18433789, 227454343, 208475153, 2204580, 98445813}))
  stage_2_butterfly_15 (
    .x_in(stage_1_per_out[30]),
    .y_in(stage_1_per_out[31]),
    .x_out(stage_2_per_in[30]),
    .y_out(stage_2_per_in[31]),
    .clk(clk),
    .rst(rst)
  );





  // TODO(Yang): stage 2 -> stage 3 permutation
  // FIXME: ignore butterfly units for now.
  stage_2_permutation #(
    .DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    .INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_2_3_per (
    .inData_0(stage_2_per_in[0]),
    .inData_1(stage_2_per_in[1]),
    .inData_2(stage_2_per_in[2]),
    .inData_3(stage_2_per_in[3]),
    .inData_4(stage_2_per_in[4]),
    .inData_5(stage_2_per_in[5]),
    .inData_6(stage_2_per_in[6]),
    .inData_7(stage_2_per_in[7]),
    .inData_8(stage_2_per_in[8]),
    .inData_9(stage_2_per_in[9]),
    .inData_10(stage_2_per_in[10]),
    .inData_11(stage_2_per_in[11]),
    .inData_12(stage_2_per_in[12]),
    .inData_13(stage_2_per_in[13]),
    .inData_14(stage_2_per_in[14]),
    .inData_15(stage_2_per_in[15]),
    .inData_16(stage_2_per_in[16]),
    .inData_17(stage_2_per_in[17]),
    .inData_18(stage_2_per_in[18]),
    .inData_19(stage_2_per_in[19]),
    .inData_20(stage_2_per_in[20]),
    .inData_21(stage_2_per_in[21]),
    .inData_22(stage_2_per_in[22]),
    .inData_23(stage_2_per_in[23]),
    .inData_24(stage_2_per_in[24]),
    .inData_25(stage_2_per_in[25]),
    .inData_26(stage_2_per_in[26]),
    .inData_27(stage_2_per_in[27]),
    .inData_28(stage_2_per_in[28]),
    .inData_29(stage_2_per_in[29]),
    .inData_30(stage_2_per_in[30]),
    .inData_31(stage_2_per_in[31]),
    .outData_0(stage_2_per_out[0]),
    .outData_1(stage_2_per_out[1]),
    .outData_2(stage_2_per_out[2]),
    .outData_3(stage_2_per_out[3]),
    .outData_4(stage_2_per_out[4]),
    .outData_5(stage_2_per_out[5]),
    .outData_6(stage_2_per_out[6]),
    .outData_7(stage_2_per_out[7]),
    .outData_8(stage_2_per_out[8]),
    .outData_9(stage_2_per_out[9]),
    .outData_10(stage_2_per_out[10]),
    .outData_11(stage_2_per_out[11]),
    .outData_12(stage_2_per_out[12]),
    .outData_13(stage_2_per_out[13]),
    .outData_14(stage_2_per_out[14]),
    .outData_15(stage_2_per_out[15]),
    .outData_16(stage_2_per_out[16]),
    .outData_17(stage_2_per_out[17]),
    .outData_18(stage_2_per_out[18]),
    .outData_19(stage_2_per_out[19]),
    .outData_20(stage_2_per_out[20]),
    .outData_21(stage_2_per_out[21]),
    .outData_22(stage_2_per_out[22]),
    .outData_23(stage_2_per_out[23]),
    .outData_24(stage_2_per_out[24]),
    .outData_25(stage_2_per_out[25]),
    .outData_26(stage_2_per_out[26]),
    .outData_27(stage_2_per_out[27]),
    .outData_28(stage_2_per_out[28]),
    .outData_29(stage_2_per_out[29]),
    .outData_30(stage_2_per_out[30]),
    .outData_31(stage_2_per_out[31]),
    .in_start(in_start[2]),
    .out_start(out_start[2]),
    .clk(clk),
    .rst(rst)
  );

  // TODO(Tian): stage 3 32 butterfly units
  butterfly #(
    .start(START_CYCLE[3]),
    .factors({135618975, 98861208, 219738759, 4839268, 141849606, 12196542, 28242170, 178386996,
              98889920, 232615475, 132483080, 102915173, 134877507, 201144768, 216395023, 167911982,
              64884498, 253800975, 42719459, 263070789, 186863562, 181295312, 168676526, 131377029,
              224068691, 205961920, 212275822, 82934386, 100123291, 23606744, 190319963, 76925614,
              209658551, 79852752, 176209504, 117274103, 99392088, 32087335, 138879618, 73081523,
              258527796, 141424302, 209725121, 68267735, 85252512, 172809179, 66242139, 68559335,
              65324949, 123440080, 49057739, 55609416, 95282463, 94612904, 262464837, 190980049,
              227819465, 181468172, 183029478, 243024363, 20857483, 16985430, 80505160, 195748297,
              198785423, 233514072, 202059197, 10720790, 1562592, 185685569, 101414187, 210770212,
              219083512, 172935357, 200399539, 236109059, 194276347, 44547301, 7460524, 222861227,
              251898247, 93740850, 34971158, 225265815, 44144526, 143102859, 103234978, 256272276,
              255286072, 109902969, 206795535, 47879495, 170930026, 164638888, 171051327, 177340471,
              224794776, 87202272, 218231468, 40718170, 176665584, 57455860, 143969870, 165350229,
              202776751, 150862394, 143779572, 43194148, 246630386, 161171966, 211426643, 200749611,
              165872957, 1613379, 247253507, 256869432, 172508742, 6010959, 242302870, 209583375,
              73698550, 225291788, 25853611, 139268485, 208297913, 215146927, 36946189, 257269778}))
  stage_3_butterfly_0 (
    .x_in(stage_2_per_out[0]),
    .y_in(stage_2_per_out[1]),
    .x_out(stage_3_per_in[0]),
    .y_out(stage_3_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({135618975, 98861208, 219738759, 4839268, 141849606, 12196542, 28242170, 178386996,
              98889920, 232615475, 132483080, 102915173, 134877507, 201144768, 216395023, 167911982,
              64884498, 253800975, 42719459, 263070789, 186863562, 181295312, 168676526, 131377029,
              224068691, 205961920, 212275822, 82934386, 100123291, 23606744, 190319963, 76925614,
              209658551, 79852752, 176209504, 117274103, 99392088, 32087335, 138879618, 73081523,
              258527796, 141424302, 209725121, 68267735, 85252512, 172809179, 66242139, 68559335,
              65324949, 123440080, 49057739, 55609416, 95282463, 94612904, 262464837, 190980049,
              227819465, 181468172, 183029478, 243024363, 20857483, 16985430, 80505160, 195748297,
              198785423, 233514072, 202059197, 10720790, 1562592, 185685569, 101414187, 210770212,
              219083512, 172935357, 200399539, 236109059, 194276347, 44547301, 7460524, 222861227,
              251898247, 93740850, 34971158, 225265815, 44144526, 143102859, 103234978, 256272276,
              255286072, 109902969, 206795535, 47879495, 170930026, 164638888, 171051327, 177340471,
              224794776, 87202272, 218231468, 40718170, 176665584, 57455860, 143969870, 165350229,
              202776751, 150862394, 143779572, 43194148, 246630386, 161171966, 211426643, 200749611,
              165872957, 1613379, 247253507, 256869432, 172508742, 6010959, 242302870, 209583375,
              73698550, 225291788, 25853611, 139268485, 208297913, 215146927, 36946189, 257269778}))
  stage_3_butterfly_1 (
    .x_in(stage_2_per_out[2]),
    .y_in(stage_2_per_out[3]),
    .x_out(stage_3_per_in[2]),
    .y_out(stage_3_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({135618975, 98861208, 219738759, 4839268, 141849606, 12196542, 28242170, 178386996,
              98889920, 232615475, 132483080, 102915173, 134877507, 201144768, 216395023, 167911982,
              64884498, 253800975, 42719459, 263070789, 186863562, 181295312, 168676526, 131377029,
              224068691, 205961920, 212275822, 82934386, 100123291, 23606744, 190319963, 76925614,
              209658551, 79852752, 176209504, 117274103, 99392088, 32087335, 138879618, 73081523,
              258527796, 141424302, 209725121, 68267735, 85252512, 172809179, 66242139, 68559335,
              65324949, 123440080, 49057739, 55609416, 95282463, 94612904, 262464837, 190980049,
              227819465, 181468172, 183029478, 243024363, 20857483, 16985430, 80505160, 195748297,
              198785423, 233514072, 202059197, 10720790, 1562592, 185685569, 101414187, 210770212,
              219083512, 172935357, 200399539, 236109059, 194276347, 44547301, 7460524, 222861227,
              251898247, 93740850, 34971158, 225265815, 44144526, 143102859, 103234978, 256272276,
              255286072, 109902969, 206795535, 47879495, 170930026, 164638888, 171051327, 177340471,
              224794776, 87202272, 218231468, 40718170, 176665584, 57455860, 143969870, 165350229,
              202776751, 150862394, 143779572, 43194148, 246630386, 161171966, 211426643, 200749611,
              165872957, 1613379, 247253507, 256869432, 172508742, 6010959, 242302870, 209583375,
              73698550, 225291788, 25853611, 139268485, 208297913, 215146927, 36946189, 257269778}))
  stage_3_butterfly_2 (
    .x_in(stage_2_per_out[4]),
    .y_in(stage_2_per_out[5]),
    .x_out(stage_3_per_in[4]),
    .y_out(stage_3_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({135618975, 98861208, 219738759, 4839268, 141849606, 12196542, 28242170, 178386996,
              98889920, 232615475, 132483080, 102915173, 134877507, 201144768, 216395023, 167911982,
              64884498, 253800975, 42719459, 263070789, 186863562, 181295312, 168676526, 131377029,
              224068691, 205961920, 212275822, 82934386, 100123291, 23606744, 190319963, 76925614,
              209658551, 79852752, 176209504, 117274103, 99392088, 32087335, 138879618, 73081523,
              258527796, 141424302, 209725121, 68267735, 85252512, 172809179, 66242139, 68559335,
              65324949, 123440080, 49057739, 55609416, 95282463, 94612904, 262464837, 190980049,
              227819465, 181468172, 183029478, 243024363, 20857483, 16985430, 80505160, 195748297,
              198785423, 233514072, 202059197, 10720790, 1562592, 185685569, 101414187, 210770212,
              219083512, 172935357, 200399539, 236109059, 194276347, 44547301, 7460524, 222861227,
              251898247, 93740850, 34971158, 225265815, 44144526, 143102859, 103234978, 256272276,
              255286072, 109902969, 206795535, 47879495, 170930026, 164638888, 171051327, 177340471,
              224794776, 87202272, 218231468, 40718170, 176665584, 57455860, 143969870, 165350229,
              202776751, 150862394, 143779572, 43194148, 246630386, 161171966, 211426643, 200749611,
              165872957, 1613379, 247253507, 256869432, 172508742, 6010959, 242302870, 209583375,
              73698550, 225291788, 25853611, 139268485, 208297913, 215146927, 36946189, 257269778}))
  stage_3_butterfly_3 (
    .x_in(stage_2_per_out[6]),
    .y_in(stage_2_per_out[7]),
    .x_out(stage_3_per_in[6]),
    .y_out(stage_3_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({135618975, 98861208, 219738759, 4839268, 141849606, 12196542, 28242170, 178386996,
              98889920, 232615475, 132483080, 102915173, 134877507, 201144768, 216395023, 167911982,
              64884498, 253800975, 42719459, 263070789, 186863562, 181295312, 168676526, 131377029,
              224068691, 205961920, 212275822, 82934386, 100123291, 23606744, 190319963, 76925614,
              209658551, 79852752, 176209504, 117274103, 99392088, 32087335, 138879618, 73081523,
              258527796, 141424302, 209725121, 68267735, 85252512, 172809179, 66242139, 68559335,
              65324949, 123440080, 49057739, 55609416, 95282463, 94612904, 262464837, 190980049,
              227819465, 181468172, 183029478, 243024363, 20857483, 16985430, 80505160, 195748297,
              198785423, 233514072, 202059197, 10720790, 1562592, 185685569, 101414187, 210770212,
              219083512, 172935357, 200399539, 236109059, 194276347, 44547301, 7460524, 222861227,
              251898247, 93740850, 34971158, 225265815, 44144526, 143102859, 103234978, 256272276,
              255286072, 109902969, 206795535, 47879495, 170930026, 164638888, 171051327, 177340471,
              224794776, 87202272, 218231468, 40718170, 176665584, 57455860, 143969870, 165350229,
              202776751, 150862394, 143779572, 43194148, 246630386, 161171966, 211426643, 200749611,
              165872957, 1613379, 247253507, 256869432, 172508742, 6010959, 242302870, 209583375,
              73698550, 225291788, 25853611, 139268485, 208297913, 215146927, 36946189, 257269778}))
  stage_3_butterfly_4 (
    .x_in(stage_2_per_out[8]),
    .y_in(stage_2_per_out[9]),
    .x_out(stage_3_per_in[8]),
    .y_out(stage_3_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({135618975, 98861208, 219738759, 4839268, 141849606, 12196542, 28242170, 178386996,
              98889920, 232615475, 132483080, 102915173, 134877507, 201144768, 216395023, 167911982,
              64884498, 253800975, 42719459, 263070789, 186863562, 181295312, 168676526, 131377029,
              224068691, 205961920, 212275822, 82934386, 100123291, 23606744, 190319963, 76925614,
              209658551, 79852752, 176209504, 117274103, 99392088, 32087335, 138879618, 73081523,
              258527796, 141424302, 209725121, 68267735, 85252512, 172809179, 66242139, 68559335,
              65324949, 123440080, 49057739, 55609416, 95282463, 94612904, 262464837, 190980049,
              227819465, 181468172, 183029478, 243024363, 20857483, 16985430, 80505160, 195748297,
              198785423, 233514072, 202059197, 10720790, 1562592, 185685569, 101414187, 210770212,
              219083512, 172935357, 200399539, 236109059, 194276347, 44547301, 7460524, 222861227,
              251898247, 93740850, 34971158, 225265815, 44144526, 143102859, 103234978, 256272276,
              255286072, 109902969, 206795535, 47879495, 170930026, 164638888, 171051327, 177340471,
              224794776, 87202272, 218231468, 40718170, 176665584, 57455860, 143969870, 165350229,
              202776751, 150862394, 143779572, 43194148, 246630386, 161171966, 211426643, 200749611,
              165872957, 1613379, 247253507, 256869432, 172508742, 6010959, 242302870, 209583375,
              73698550, 225291788, 25853611, 139268485, 208297913, 215146927, 36946189, 257269778}))
  stage_3_butterfly_5 (
    .x_in(stage_2_per_out[10]),
    .y_in(stage_2_per_out[11]),
    .x_out(stage_3_per_in[10]),
    .y_out(stage_3_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({135618975, 98861208, 219738759, 4839268, 141849606, 12196542, 28242170, 178386996,
              98889920, 232615475, 132483080, 102915173, 134877507, 201144768, 216395023, 167911982,
              64884498, 253800975, 42719459, 263070789, 186863562, 181295312, 168676526, 131377029,
              224068691, 205961920, 212275822, 82934386, 100123291, 23606744, 190319963, 76925614,
              209658551, 79852752, 176209504, 117274103, 99392088, 32087335, 138879618, 73081523,
              258527796, 141424302, 209725121, 68267735, 85252512, 172809179, 66242139, 68559335,
              65324949, 123440080, 49057739, 55609416, 95282463, 94612904, 262464837, 190980049,
              227819465, 181468172, 183029478, 243024363, 20857483, 16985430, 80505160, 195748297,
              198785423, 233514072, 202059197, 10720790, 1562592, 185685569, 101414187, 210770212,
              219083512, 172935357, 200399539, 236109059, 194276347, 44547301, 7460524, 222861227,
              251898247, 93740850, 34971158, 225265815, 44144526, 143102859, 103234978, 256272276,
              255286072, 109902969, 206795535, 47879495, 170930026, 164638888, 171051327, 177340471,
              224794776, 87202272, 218231468, 40718170, 176665584, 57455860, 143969870, 165350229,
              202776751, 150862394, 143779572, 43194148, 246630386, 161171966, 211426643, 200749611,
              165872957, 1613379, 247253507, 256869432, 172508742, 6010959, 242302870, 209583375,
              73698550, 225291788, 25853611, 139268485, 208297913, 215146927, 36946189, 257269778}))
  stage_3_butterfly_6 (
    .x_in(stage_2_per_out[12]),
    .y_in(stage_2_per_out[13]),
    .x_out(stage_3_per_in[12]),
    .y_out(stage_3_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({135618975, 98861208, 219738759, 4839268, 141849606, 12196542, 28242170, 178386996,
              98889920, 232615475, 132483080, 102915173, 134877507, 201144768, 216395023, 167911982,
              64884498, 253800975, 42719459, 263070789, 186863562, 181295312, 168676526, 131377029,
              224068691, 205961920, 212275822, 82934386, 100123291, 23606744, 190319963, 76925614,
              209658551, 79852752, 176209504, 117274103, 99392088, 32087335, 138879618, 73081523,
              258527796, 141424302, 209725121, 68267735, 85252512, 172809179, 66242139, 68559335,
              65324949, 123440080, 49057739, 55609416, 95282463, 94612904, 262464837, 190980049,
              227819465, 181468172, 183029478, 243024363, 20857483, 16985430, 80505160, 195748297,
              198785423, 233514072, 202059197, 10720790, 1562592, 185685569, 101414187, 210770212,
              219083512, 172935357, 200399539, 236109059, 194276347, 44547301, 7460524, 222861227,
              251898247, 93740850, 34971158, 225265815, 44144526, 143102859, 103234978, 256272276,
              255286072, 109902969, 206795535, 47879495, 170930026, 164638888, 171051327, 177340471,
              224794776, 87202272, 218231468, 40718170, 176665584, 57455860, 143969870, 165350229,
              202776751, 150862394, 143779572, 43194148, 246630386, 161171966, 211426643, 200749611,
              165872957, 1613379, 247253507, 256869432, 172508742, 6010959, 242302870, 209583375,
              73698550, 225291788, 25853611, 139268485, 208297913, 215146927, 36946189, 257269778}))
  stage_3_butterfly_7 (
    .x_in(stage_2_per_out[14]),
    .y_in(stage_2_per_out[15]),
    .x_out(stage_3_per_in[14]),
    .y_out(stage_3_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({42355602, 77981460, 24688427, 233888407, 45686070, 199633043, 110403916, 23405380,
              78649100, 142181410, 170284131, 169182486, 17861009, 160841949, 202071175, 254132077,
              160254284, 8411857, 224586596, 34256894, 57574719, 100229847, 181281889, 79136411,
              117221766, 75073484, 205290416, 109479656, 182702557, 13458851, 65413984, 205525433,
              136878682, 192832423, 129576773, 60548134, 5829490, 56246211, 61644903, 140366124,
              61345534, 62117518, 263077695, 210734246, 148801771, 148390399, 67321994, 149992379,
              69773246, 209085090, 196771169, 50986641, 56155754, 10003248, 82155735, 114486793,
              137065607, 241313184, 155060883, 266671862, 40158424, 25944135, 207329882, 184310992,
              54534442, 212802310, 258226806, 237102043, 249146534, 50222736, 219898221, 131023241,
              61720173, 18298478, 167366585, 229100654, 64764693, 209886001, 93469550, 196522490,
              258559590, 145034471, 68493159, 185138250, 134269022, 186841927, 63483304, 122332647,
              184644727, 160807241, 225389748, 247289727, 142306631, 258257144, 95251863, 196328787,
              220994759, 193915204, 17231623, 154421517, 8950678, 92650808, 252241817, 238382196,
              225784463, 171362072, 156366160, 171541778, 61664240, 30930936, 35918322, 61997323,
              23892097, 158727274, 35924353, 242025902, 234350511, 226213489, 6574921, 137672988,
              49504466, 244216783, 119169851, 49675259, 66505970, 158168844, 6292910, 182691070}))
  stage_3_butterfly_8 (
    .x_in(stage_2_per_out[16]),
    .y_in(stage_2_per_out[17]),
    .x_out(stage_3_per_in[16]),
    .y_out(stage_3_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({42355602, 77981460, 24688427, 233888407, 45686070, 199633043, 110403916, 23405380,
              78649100, 142181410, 170284131, 169182486, 17861009, 160841949, 202071175, 254132077,
              160254284, 8411857, 224586596, 34256894, 57574719, 100229847, 181281889, 79136411,
              117221766, 75073484, 205290416, 109479656, 182702557, 13458851, 65413984, 205525433,
              136878682, 192832423, 129576773, 60548134, 5829490, 56246211, 61644903, 140366124,
              61345534, 62117518, 263077695, 210734246, 148801771, 148390399, 67321994, 149992379,
              69773246, 209085090, 196771169, 50986641, 56155754, 10003248, 82155735, 114486793,
              137065607, 241313184, 155060883, 266671862, 40158424, 25944135, 207329882, 184310992,
              54534442, 212802310, 258226806, 237102043, 249146534, 50222736, 219898221, 131023241,
              61720173, 18298478, 167366585, 229100654, 64764693, 209886001, 93469550, 196522490,
              258559590, 145034471, 68493159, 185138250, 134269022, 186841927, 63483304, 122332647,
              184644727, 160807241, 225389748, 247289727, 142306631, 258257144, 95251863, 196328787,
              220994759, 193915204, 17231623, 154421517, 8950678, 92650808, 252241817, 238382196,
              225784463, 171362072, 156366160, 171541778, 61664240, 30930936, 35918322, 61997323,
              23892097, 158727274, 35924353, 242025902, 234350511, 226213489, 6574921, 137672988,
              49504466, 244216783, 119169851, 49675259, 66505970, 158168844, 6292910, 182691070}))
  stage_3_butterfly_9 (
    .x_in(stage_2_per_out[18]),
    .y_in(stage_2_per_out[19]),
    .x_out(stage_3_per_in[18]),
    .y_out(stage_3_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({42355602, 77981460, 24688427, 233888407, 45686070, 199633043, 110403916, 23405380,
              78649100, 142181410, 170284131, 169182486, 17861009, 160841949, 202071175, 254132077,
              160254284, 8411857, 224586596, 34256894, 57574719, 100229847, 181281889, 79136411,
              117221766, 75073484, 205290416, 109479656, 182702557, 13458851, 65413984, 205525433,
              136878682, 192832423, 129576773, 60548134, 5829490, 56246211, 61644903, 140366124,
              61345534, 62117518, 263077695, 210734246, 148801771, 148390399, 67321994, 149992379,
              69773246, 209085090, 196771169, 50986641, 56155754, 10003248, 82155735, 114486793,
              137065607, 241313184, 155060883, 266671862, 40158424, 25944135, 207329882, 184310992,
              54534442, 212802310, 258226806, 237102043, 249146534, 50222736, 219898221, 131023241,
              61720173, 18298478, 167366585, 229100654, 64764693, 209886001, 93469550, 196522490,
              258559590, 145034471, 68493159, 185138250, 134269022, 186841927, 63483304, 122332647,
              184644727, 160807241, 225389748, 247289727, 142306631, 258257144, 95251863, 196328787,
              220994759, 193915204, 17231623, 154421517, 8950678, 92650808, 252241817, 238382196,
              225784463, 171362072, 156366160, 171541778, 61664240, 30930936, 35918322, 61997323,
              23892097, 158727274, 35924353, 242025902, 234350511, 226213489, 6574921, 137672988,
              49504466, 244216783, 119169851, 49675259, 66505970, 158168844, 6292910, 182691070}))
  stage_3_butterfly_10 (
    .x_in(stage_2_per_out[20]),
    .y_in(stage_2_per_out[21]),
    .x_out(stage_3_per_in[20]),
    .y_out(stage_3_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({42355602, 77981460, 24688427, 233888407, 45686070, 199633043, 110403916, 23405380,
              78649100, 142181410, 170284131, 169182486, 17861009, 160841949, 202071175, 254132077,
              160254284, 8411857, 224586596, 34256894, 57574719, 100229847, 181281889, 79136411,
              117221766, 75073484, 205290416, 109479656, 182702557, 13458851, 65413984, 205525433,
              136878682, 192832423, 129576773, 60548134, 5829490, 56246211, 61644903, 140366124,
              61345534, 62117518, 263077695, 210734246, 148801771, 148390399, 67321994, 149992379,
              69773246, 209085090, 196771169, 50986641, 56155754, 10003248, 82155735, 114486793,
              137065607, 241313184, 155060883, 266671862, 40158424, 25944135, 207329882, 184310992,
              54534442, 212802310, 258226806, 237102043, 249146534, 50222736, 219898221, 131023241,
              61720173, 18298478, 167366585, 229100654, 64764693, 209886001, 93469550, 196522490,
              258559590, 145034471, 68493159, 185138250, 134269022, 186841927, 63483304, 122332647,
              184644727, 160807241, 225389748, 247289727, 142306631, 258257144, 95251863, 196328787,
              220994759, 193915204, 17231623, 154421517, 8950678, 92650808, 252241817, 238382196,
              225784463, 171362072, 156366160, 171541778, 61664240, 30930936, 35918322, 61997323,
              23892097, 158727274, 35924353, 242025902, 234350511, 226213489, 6574921, 137672988,
              49504466, 244216783, 119169851, 49675259, 66505970, 158168844, 6292910, 182691070}))
  stage_3_butterfly_11 (
    .x_in(stage_2_per_out[22]),
    .y_in(stage_2_per_out[23]),
    .x_out(stage_3_per_in[22]),
    .y_out(stage_3_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({42355602, 77981460, 24688427, 233888407, 45686070, 199633043, 110403916, 23405380,
              78649100, 142181410, 170284131, 169182486, 17861009, 160841949, 202071175, 254132077,
              160254284, 8411857, 224586596, 34256894, 57574719, 100229847, 181281889, 79136411,
              117221766, 75073484, 205290416, 109479656, 182702557, 13458851, 65413984, 205525433,
              136878682, 192832423, 129576773, 60548134, 5829490, 56246211, 61644903, 140366124,
              61345534, 62117518, 263077695, 210734246, 148801771, 148390399, 67321994, 149992379,
              69773246, 209085090, 196771169, 50986641, 56155754, 10003248, 82155735, 114486793,
              137065607, 241313184, 155060883, 266671862, 40158424, 25944135, 207329882, 184310992,
              54534442, 212802310, 258226806, 237102043, 249146534, 50222736, 219898221, 131023241,
              61720173, 18298478, 167366585, 229100654, 64764693, 209886001, 93469550, 196522490,
              258559590, 145034471, 68493159, 185138250, 134269022, 186841927, 63483304, 122332647,
              184644727, 160807241, 225389748, 247289727, 142306631, 258257144, 95251863, 196328787,
              220994759, 193915204, 17231623, 154421517, 8950678, 92650808, 252241817, 238382196,
              225784463, 171362072, 156366160, 171541778, 61664240, 30930936, 35918322, 61997323,
              23892097, 158727274, 35924353, 242025902, 234350511, 226213489, 6574921, 137672988,
              49504466, 244216783, 119169851, 49675259, 66505970, 158168844, 6292910, 182691070}))
  stage_3_butterfly_12 (
    .x_in(stage_2_per_out[24]),
    .y_in(stage_2_per_out[25]),
    .x_out(stage_3_per_in[24]),
    .y_out(stage_3_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({42355602, 77981460, 24688427, 233888407, 45686070, 199633043, 110403916, 23405380,
              78649100, 142181410, 170284131, 169182486, 17861009, 160841949, 202071175, 254132077,
              160254284, 8411857, 224586596, 34256894, 57574719, 100229847, 181281889, 79136411,
              117221766, 75073484, 205290416, 109479656, 182702557, 13458851, 65413984, 205525433,
              136878682, 192832423, 129576773, 60548134, 5829490, 56246211, 61644903, 140366124,
              61345534, 62117518, 263077695, 210734246, 148801771, 148390399, 67321994, 149992379,
              69773246, 209085090, 196771169, 50986641, 56155754, 10003248, 82155735, 114486793,
              137065607, 241313184, 155060883, 266671862, 40158424, 25944135, 207329882, 184310992,
              54534442, 212802310, 258226806, 237102043, 249146534, 50222736, 219898221, 131023241,
              61720173, 18298478, 167366585, 229100654, 64764693, 209886001, 93469550, 196522490,
              258559590, 145034471, 68493159, 185138250, 134269022, 186841927, 63483304, 122332647,
              184644727, 160807241, 225389748, 247289727, 142306631, 258257144, 95251863, 196328787,
              220994759, 193915204, 17231623, 154421517, 8950678, 92650808, 252241817, 238382196,
              225784463, 171362072, 156366160, 171541778, 61664240, 30930936, 35918322, 61997323,
              23892097, 158727274, 35924353, 242025902, 234350511, 226213489, 6574921, 137672988,
              49504466, 244216783, 119169851, 49675259, 66505970, 158168844, 6292910, 182691070}))
  stage_3_butterfly_13 (
    .x_in(stage_2_per_out[26]),
    .y_in(stage_2_per_out[27]),
    .x_out(stage_3_per_in[26]),
    .y_out(stage_3_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({42355602, 77981460, 24688427, 233888407, 45686070, 199633043, 110403916, 23405380,
              78649100, 142181410, 170284131, 169182486, 17861009, 160841949, 202071175, 254132077,
              160254284, 8411857, 224586596, 34256894, 57574719, 100229847, 181281889, 79136411,
              117221766, 75073484, 205290416, 109479656, 182702557, 13458851, 65413984, 205525433,
              136878682, 192832423, 129576773, 60548134, 5829490, 56246211, 61644903, 140366124,
              61345534, 62117518, 263077695, 210734246, 148801771, 148390399, 67321994, 149992379,
              69773246, 209085090, 196771169, 50986641, 56155754, 10003248, 82155735, 114486793,
              137065607, 241313184, 155060883, 266671862, 40158424, 25944135, 207329882, 184310992,
              54534442, 212802310, 258226806, 237102043, 249146534, 50222736, 219898221, 131023241,
              61720173, 18298478, 167366585, 229100654, 64764693, 209886001, 93469550, 196522490,
              258559590, 145034471, 68493159, 185138250, 134269022, 186841927, 63483304, 122332647,
              184644727, 160807241, 225389748, 247289727, 142306631, 258257144, 95251863, 196328787,
              220994759, 193915204, 17231623, 154421517, 8950678, 92650808, 252241817, 238382196,
              225784463, 171362072, 156366160, 171541778, 61664240, 30930936, 35918322, 61997323,
              23892097, 158727274, 35924353, 242025902, 234350511, 226213489, 6574921, 137672988,
              49504466, 244216783, 119169851, 49675259, 66505970, 158168844, 6292910, 182691070}))
  stage_3_butterfly_14 (
    .x_in(stage_2_per_out[28]),
    .y_in(stage_2_per_out[29]),
    .x_out(stage_3_per_in[28]),
    .y_out(stage_3_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[3]),
    .factors({42355602, 77981460, 24688427, 233888407, 45686070, 199633043, 110403916, 23405380,
              78649100, 142181410, 170284131, 169182486, 17861009, 160841949, 202071175, 254132077,
              160254284, 8411857, 224586596, 34256894, 57574719, 100229847, 181281889, 79136411,
              117221766, 75073484, 205290416, 109479656, 182702557, 13458851, 65413984, 205525433,
              136878682, 192832423, 129576773, 60548134, 5829490, 56246211, 61644903, 140366124,
              61345534, 62117518, 263077695, 210734246, 148801771, 148390399, 67321994, 149992379,
              69773246, 209085090, 196771169, 50986641, 56155754, 10003248, 82155735, 114486793,
              137065607, 241313184, 155060883, 266671862, 40158424, 25944135, 207329882, 184310992,
              54534442, 212802310, 258226806, 237102043, 249146534, 50222736, 219898221, 131023241,
              61720173, 18298478, 167366585, 229100654, 64764693, 209886001, 93469550, 196522490,
              258559590, 145034471, 68493159, 185138250, 134269022, 186841927, 63483304, 122332647,
              184644727, 160807241, 225389748, 247289727, 142306631, 258257144, 95251863, 196328787,
              220994759, 193915204, 17231623, 154421517, 8950678, 92650808, 252241817, 238382196,
              225784463, 171362072, 156366160, 171541778, 61664240, 30930936, 35918322, 61997323,
              23892097, 158727274, 35924353, 242025902, 234350511, 226213489, 6574921, 137672988,
              49504466, 244216783, 119169851, 49675259, 66505970, 158168844, 6292910, 182691070}))
  stage_3_butterfly_15 (
    .x_in(stage_2_per_out[30]),
    .y_in(stage_2_per_out[31]),
    .x_out(stage_3_per_in[30]),
    .y_out(stage_3_per_in[31]),
    .clk(clk),
    .rst(rst)
  );




  // TODO(Yang): stage 3 -> stage 4 permutation
  // FIXME: ignore butterfly units for now.
  stage_3_permutation #(
    .DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    .INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_3_4_per (
    .inData_0(stage_3_per_in[0]),
    .inData_1(stage_3_per_in[1]),
    .inData_2(stage_3_per_in[2]),
    .inData_3(stage_3_per_in[3]),
    .inData_4(stage_3_per_in[4]),
    .inData_5(stage_3_per_in[5]),
    .inData_6(stage_3_per_in[6]),
    .inData_7(stage_3_per_in[7]),
    .inData_8(stage_3_per_in[8]),
    .inData_9(stage_3_per_in[9]),
    .inData_10(stage_3_per_in[10]),
    .inData_11(stage_3_per_in[11]),
    .inData_12(stage_3_per_in[12]),
    .inData_13(stage_3_per_in[13]),
    .inData_14(stage_3_per_in[14]),
    .inData_15(stage_3_per_in[15]),
    .inData_16(stage_3_per_in[16]),
    .inData_17(stage_3_per_in[17]),
    .inData_18(stage_3_per_in[18]),
    .inData_19(stage_3_per_in[19]),
    .inData_20(stage_3_per_in[20]),
    .inData_21(stage_3_per_in[21]),
    .inData_22(stage_3_per_in[22]),
    .inData_23(stage_3_per_in[23]),
    .inData_24(stage_3_per_in[24]),
    .inData_25(stage_3_per_in[25]),
    .inData_26(stage_3_per_in[26]),
    .inData_27(stage_3_per_in[27]),
    .inData_28(stage_3_per_in[28]),
    .inData_29(stage_3_per_in[29]),
    .inData_30(stage_3_per_in[30]),
    .inData_31(stage_3_per_in[31]),
    .outData_0(stage_3_per_out[0]),
    .outData_1(stage_3_per_out[1]),
    .outData_2(stage_3_per_out[2]),
    .outData_3(stage_3_per_out[3]),
    .outData_4(stage_3_per_out[4]),
    .outData_5(stage_3_per_out[5]),
    .outData_6(stage_3_per_out[6]),
    .outData_7(stage_3_per_out[7]),
    .outData_8(stage_3_per_out[8]),
    .outData_9(stage_3_per_out[9]),
    .outData_10(stage_3_per_out[10]),
    .outData_11(stage_3_per_out[11]),
    .outData_12(stage_3_per_out[12]),
    .outData_13(stage_3_per_out[13]),
    .outData_14(stage_3_per_out[14]),
    .outData_15(stage_3_per_out[15]),
    .outData_16(stage_3_per_out[16]),
    .outData_17(stage_3_per_out[17]),
    .outData_18(stage_3_per_out[18]),
    .outData_19(stage_3_per_out[19]),
    .outData_20(stage_3_per_out[20]),
    .outData_21(stage_3_per_out[21]),
    .outData_22(stage_3_per_out[22]),
    .outData_23(stage_3_per_out[23]),
    .outData_24(stage_3_per_out[24]),
    .outData_25(stage_3_per_out[25]),
    .outData_26(stage_3_per_out[26]),
    .outData_27(stage_3_per_out[27]),
    .outData_28(stage_3_per_out[28]),
    .outData_29(stage_3_per_out[29]),
    .outData_30(stage_3_per_out[30]),
    .outData_31(stage_3_per_out[31]),
    .in_start(in_start[3]),
    .out_start(out_start[3]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 4 32 butterfly units
  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 261793746, 116401819, 18729522, 11101448, 68136911, 71064168, 166886297,
              189762285, 21713495, 81956368, 176917280, 244883276, 7055647, 135288005, 238498066,
              229228230, 148662095, 216143425, 181639510, 101839787, 256040960, 265950570, 240677074,
              85922744, 123185272, 254450415, 97765534, 10571783, 170227406, 14542514, 40475021,
              117496916, 193371292, 250166212, 167885779, 192696288, 159404461, 130557622, 37051834,
              106640438, 183348420, 234030247, 41155851, 90597117, 173702965, 209086118, 258612781,
              189881206, 186592442, 10130658, 139182289, 241125460, 243304319, 176471684, 83853696,
              209161759, 236144340, 231358848, 230433664, 245906264, 189591954, 63350037, 54284329,
              55721255, 254509489, 47751177, 15417588, 64217206, 66148505, 229216409, 108083129,
              40553702, 118518376, 204666342, 241682233, 214551729, 108810259, 33479018, 223427563,
              226739459, 67012048, 34119889, 77337691, 246744565, 104174682, 2795054, 161827885,
              104557084, 155168409, 96142103, 118841873, 104784816, 3883583, 41086336, 134866823,
              122008382, 25569479, 211668928, 123954975, 225636920, 120936039, 197074908, 210298252,
              47994339, 13519489, 252442032, 162031725, 168407516, 132703565, 9720223, 19493867,
              184226747, 71933862, 143969713, 230702770, 69161747, 180525688, 245828202, 13250338,
              239545014, 139555205, 98878775, 9446767, 72738487, 171721518, 217644581, 249970613}))
  stage_4_butterfly_0 (
    .x_in(stage_3_per_out[0]),
    .y_in(stage_3_per_out[1]),
    .x_out(stage_4_per_in[0]),
    .y_out(stage_4_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 261793746, 116401819, 18729522, 11101448, 68136911, 71064168, 166886297,
              189762285, 21713495, 81956368, 176917280, 244883276, 7055647, 135288005, 238498066,
              229228230, 148662095, 216143425, 181639510, 101839787, 256040960, 265950570, 240677074,
              85922744, 123185272, 254450415, 97765534, 10571783, 170227406, 14542514, 40475021,
              117496916, 193371292, 250166212, 167885779, 192696288, 159404461, 130557622, 37051834,
              106640438, 183348420, 234030247, 41155851, 90597117, 173702965, 209086118, 258612781,
              189881206, 186592442, 10130658, 139182289, 241125460, 243304319, 176471684, 83853696,
              209161759, 236144340, 231358848, 230433664, 245906264, 189591954, 63350037, 54284329,
              55721255, 254509489, 47751177, 15417588, 64217206, 66148505, 229216409, 108083129,
              40553702, 118518376, 204666342, 241682233, 214551729, 108810259, 33479018, 223427563,
              226739459, 67012048, 34119889, 77337691, 246744565, 104174682, 2795054, 161827885,
              104557084, 155168409, 96142103, 118841873, 104784816, 3883583, 41086336, 134866823,
              122008382, 25569479, 211668928, 123954975, 225636920, 120936039, 197074908, 210298252,
              47994339, 13519489, 252442032, 162031725, 168407516, 132703565, 9720223, 19493867,
              184226747, 71933862, 143969713, 230702770, 69161747, 180525688, 245828202, 13250338,
              239545014, 139555205, 98878775, 9446767, 72738487, 171721518, 217644581, 249970613}))
  stage_4_butterfly_1 (
    .x_in(stage_3_per_out[2]),
    .y_in(stage_3_per_out[3]),
    .x_out(stage_4_per_in[2]),
    .y_out(stage_4_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 261793746, 116401819, 18729522, 11101448, 68136911, 71064168, 166886297,
              189762285, 21713495, 81956368, 176917280, 244883276, 7055647, 135288005, 238498066,
              229228230, 148662095, 216143425, 181639510, 101839787, 256040960, 265950570, 240677074,
              85922744, 123185272, 254450415, 97765534, 10571783, 170227406, 14542514, 40475021,
              117496916, 193371292, 250166212, 167885779, 192696288, 159404461, 130557622, 37051834,
              106640438, 183348420, 234030247, 41155851, 90597117, 173702965, 209086118, 258612781,
              189881206, 186592442, 10130658, 139182289, 241125460, 243304319, 176471684, 83853696,
              209161759, 236144340, 231358848, 230433664, 245906264, 189591954, 63350037, 54284329,
              55721255, 254509489, 47751177, 15417588, 64217206, 66148505, 229216409, 108083129,
              40553702, 118518376, 204666342, 241682233, 214551729, 108810259, 33479018, 223427563,
              226739459, 67012048, 34119889, 77337691, 246744565, 104174682, 2795054, 161827885,
              104557084, 155168409, 96142103, 118841873, 104784816, 3883583, 41086336, 134866823,
              122008382, 25569479, 211668928, 123954975, 225636920, 120936039, 197074908, 210298252,
              47994339, 13519489, 252442032, 162031725, 168407516, 132703565, 9720223, 19493867,
              184226747, 71933862, 143969713, 230702770, 69161747, 180525688, 245828202, 13250338,
              239545014, 139555205, 98878775, 9446767, 72738487, 171721518, 217644581, 249970613}))
  stage_4_butterfly_2 (
    .x_in(stage_3_per_out[4]),
    .y_in(stage_3_per_out[5]),
    .x_out(stage_4_per_in[4]),
    .y_out(stage_4_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 261793746, 116401819, 18729522, 11101448, 68136911, 71064168, 166886297,
              189762285, 21713495, 81956368, 176917280, 244883276, 7055647, 135288005, 238498066,
              229228230, 148662095, 216143425, 181639510, 101839787, 256040960, 265950570, 240677074,
              85922744, 123185272, 254450415, 97765534, 10571783, 170227406, 14542514, 40475021,
              117496916, 193371292, 250166212, 167885779, 192696288, 159404461, 130557622, 37051834,
              106640438, 183348420, 234030247, 41155851, 90597117, 173702965, 209086118, 258612781,
              189881206, 186592442, 10130658, 139182289, 241125460, 243304319, 176471684, 83853696,
              209161759, 236144340, 231358848, 230433664, 245906264, 189591954, 63350037, 54284329,
              55721255, 254509489, 47751177, 15417588, 64217206, 66148505, 229216409, 108083129,
              40553702, 118518376, 204666342, 241682233, 214551729, 108810259, 33479018, 223427563,
              226739459, 67012048, 34119889, 77337691, 246744565, 104174682, 2795054, 161827885,
              104557084, 155168409, 96142103, 118841873, 104784816, 3883583, 41086336, 134866823,
              122008382, 25569479, 211668928, 123954975, 225636920, 120936039, 197074908, 210298252,
              47994339, 13519489, 252442032, 162031725, 168407516, 132703565, 9720223, 19493867,
              184226747, 71933862, 143969713, 230702770, 69161747, 180525688, 245828202, 13250338,
              239545014, 139555205, 98878775, 9446767, 72738487, 171721518, 217644581, 249970613}))
  stage_4_butterfly_3 (
    .x_in(stage_3_per_out[6]),
    .y_in(stage_3_per_out[7]),
    .x_out(stage_4_per_in[6]),
    .y_out(stage_4_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 261793746, 116401819, 18729522, 11101448, 68136911, 71064168, 166886297,
              189762285, 21713495, 81956368, 176917280, 244883276, 7055647, 135288005, 238498066,
              229228230, 148662095, 216143425, 181639510, 101839787, 256040960, 265950570, 240677074,
              85922744, 123185272, 254450415, 97765534, 10571783, 170227406, 14542514, 40475021,
              117496916, 193371292, 250166212, 167885779, 192696288, 159404461, 130557622, 37051834,
              106640438, 183348420, 234030247, 41155851, 90597117, 173702965, 209086118, 258612781,
              189881206, 186592442, 10130658, 139182289, 241125460, 243304319, 176471684, 83853696,
              209161759, 236144340, 231358848, 230433664, 245906264, 189591954, 63350037, 54284329,
              55721255, 254509489, 47751177, 15417588, 64217206, 66148505, 229216409, 108083129,
              40553702, 118518376, 204666342, 241682233, 214551729, 108810259, 33479018, 223427563,
              226739459, 67012048, 34119889, 77337691, 246744565, 104174682, 2795054, 161827885,
              104557084, 155168409, 96142103, 118841873, 104784816, 3883583, 41086336, 134866823,
              122008382, 25569479, 211668928, 123954975, 225636920, 120936039, 197074908, 210298252,
              47994339, 13519489, 252442032, 162031725, 168407516, 132703565, 9720223, 19493867,
              184226747, 71933862, 143969713, 230702770, 69161747, 180525688, 245828202, 13250338,
              239545014, 139555205, 98878775, 9446767, 72738487, 171721518, 217644581, 249970613}))
  stage_4_butterfly_4 (
    .x_in(stage_3_per_out[8]),
    .y_in(stage_3_per_out[9]),
    .x_out(stage_4_per_in[8]),
    .y_out(stage_4_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 261793746, 116401819, 18729522, 11101448, 68136911, 71064168, 166886297,
              189762285, 21713495, 81956368, 176917280, 244883276, 7055647, 135288005, 238498066,
              229228230, 148662095, 216143425, 181639510, 101839787, 256040960, 265950570, 240677074,
              85922744, 123185272, 254450415, 97765534, 10571783, 170227406, 14542514, 40475021,
              117496916, 193371292, 250166212, 167885779, 192696288, 159404461, 130557622, 37051834,
              106640438, 183348420, 234030247, 41155851, 90597117, 173702965, 209086118, 258612781,
              189881206, 186592442, 10130658, 139182289, 241125460, 243304319, 176471684, 83853696,
              209161759, 236144340, 231358848, 230433664, 245906264, 189591954, 63350037, 54284329,
              55721255, 254509489, 47751177, 15417588, 64217206, 66148505, 229216409, 108083129,
              40553702, 118518376, 204666342, 241682233, 214551729, 108810259, 33479018, 223427563,
              226739459, 67012048, 34119889, 77337691, 246744565, 104174682, 2795054, 161827885,
              104557084, 155168409, 96142103, 118841873, 104784816, 3883583, 41086336, 134866823,
              122008382, 25569479, 211668928, 123954975, 225636920, 120936039, 197074908, 210298252,
              47994339, 13519489, 252442032, 162031725, 168407516, 132703565, 9720223, 19493867,
              184226747, 71933862, 143969713, 230702770, 69161747, 180525688, 245828202, 13250338,
              239545014, 139555205, 98878775, 9446767, 72738487, 171721518, 217644581, 249970613}))
  stage_4_butterfly_5 (
    .x_in(stage_3_per_out[10]),
    .y_in(stage_3_per_out[11]),
    .x_out(stage_4_per_in[10]),
    .y_out(stage_4_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 261793746, 116401819, 18729522, 11101448, 68136911, 71064168, 166886297,
              189762285, 21713495, 81956368, 176917280, 244883276, 7055647, 135288005, 238498066,
              229228230, 148662095, 216143425, 181639510, 101839787, 256040960, 265950570, 240677074,
              85922744, 123185272, 254450415, 97765534, 10571783, 170227406, 14542514, 40475021,
              117496916, 193371292, 250166212, 167885779, 192696288, 159404461, 130557622, 37051834,
              106640438, 183348420, 234030247, 41155851, 90597117, 173702965, 209086118, 258612781,
              189881206, 186592442, 10130658, 139182289, 241125460, 243304319, 176471684, 83853696,
              209161759, 236144340, 231358848, 230433664, 245906264, 189591954, 63350037, 54284329,
              55721255, 254509489, 47751177, 15417588, 64217206, 66148505, 229216409, 108083129,
              40553702, 118518376, 204666342, 241682233, 214551729, 108810259, 33479018, 223427563,
              226739459, 67012048, 34119889, 77337691, 246744565, 104174682, 2795054, 161827885,
              104557084, 155168409, 96142103, 118841873, 104784816, 3883583, 41086336, 134866823,
              122008382, 25569479, 211668928, 123954975, 225636920, 120936039, 197074908, 210298252,
              47994339, 13519489, 252442032, 162031725, 168407516, 132703565, 9720223, 19493867,
              184226747, 71933862, 143969713, 230702770, 69161747, 180525688, 245828202, 13250338,
              239545014, 139555205, 98878775, 9446767, 72738487, 171721518, 217644581, 249970613}))
  stage_4_butterfly_6 (
    .x_in(stage_3_per_out[12]),
    .y_in(stage_3_per_out[13]),
    .x_out(stage_4_per_in[12]),
    .y_out(stage_4_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 261793746, 116401819, 18729522, 11101448, 68136911, 71064168, 166886297,
              189762285, 21713495, 81956368, 176917280, 244883276, 7055647, 135288005, 238498066,
              229228230, 148662095, 216143425, 181639510, 101839787, 256040960, 265950570, 240677074,
              85922744, 123185272, 254450415, 97765534, 10571783, 170227406, 14542514, 40475021,
              117496916, 193371292, 250166212, 167885779, 192696288, 159404461, 130557622, 37051834,
              106640438, 183348420, 234030247, 41155851, 90597117, 173702965, 209086118, 258612781,
              189881206, 186592442, 10130658, 139182289, 241125460, 243304319, 176471684, 83853696,
              209161759, 236144340, 231358848, 230433664, 245906264, 189591954, 63350037, 54284329,
              55721255, 254509489, 47751177, 15417588, 64217206, 66148505, 229216409, 108083129,
              40553702, 118518376, 204666342, 241682233, 214551729, 108810259, 33479018, 223427563,
              226739459, 67012048, 34119889, 77337691, 246744565, 104174682, 2795054, 161827885,
              104557084, 155168409, 96142103, 118841873, 104784816, 3883583, 41086336, 134866823,
              122008382, 25569479, 211668928, 123954975, 225636920, 120936039, 197074908, 210298252,
              47994339, 13519489, 252442032, 162031725, 168407516, 132703565, 9720223, 19493867,
              184226747, 71933862, 143969713, 230702770, 69161747, 180525688, 245828202, 13250338,
              239545014, 139555205, 98878775, 9446767, 72738487, 171721518, 217644581, 249970613}))
  stage_4_butterfly_7 (
    .x_in(stage_3_per_out[14]),
    .y_in(stage_3_per_out[15]),
    .x_out(stage_4_per_in[14]),
    .y_out(stage_4_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 261793746, 116401819, 18729522, 11101448, 68136911, 71064168, 166886297,
              189762285, 21713495, 81956368, 176917280, 244883276, 7055647, 135288005, 238498066,
              229228230, 148662095, 216143425, 181639510, 101839787, 256040960, 265950570, 240677074,
              85922744, 123185272, 254450415, 97765534, 10571783, 170227406, 14542514, 40475021,
              117496916, 193371292, 250166212, 167885779, 192696288, 159404461, 130557622, 37051834,
              106640438, 183348420, 234030247, 41155851, 90597117, 173702965, 209086118, 258612781,
              189881206, 186592442, 10130658, 139182289, 241125460, 243304319, 176471684, 83853696,
              209161759, 236144340, 231358848, 230433664, 245906264, 189591954, 63350037, 54284329,
              55721255, 254509489, 47751177, 15417588, 64217206, 66148505, 229216409, 108083129,
              40553702, 118518376, 204666342, 241682233, 214551729, 108810259, 33479018, 223427563,
              226739459, 67012048, 34119889, 77337691, 246744565, 104174682, 2795054, 161827885,
              104557084, 155168409, 96142103, 118841873, 104784816, 3883583, 41086336, 134866823,
              122008382, 25569479, 211668928, 123954975, 225636920, 120936039, 197074908, 210298252,
              47994339, 13519489, 252442032, 162031725, 168407516, 132703565, 9720223, 19493867,
              184226747, 71933862, 143969713, 230702770, 69161747, 180525688, 245828202, 13250338,
              239545014, 139555205, 98878775, 9446767, 72738487, 171721518, 217644581, 249970613}))
  stage_4_butterfly_8 (
    .x_in(stage_3_per_out[16]),
    .y_in(stage_3_per_out[17]),
    .x_out(stage_4_per_in[16]),
    .y_out(stage_4_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 261793746, 116401819, 18729522, 11101448, 68136911, 71064168, 166886297,
              189762285, 21713495, 81956368, 176917280, 244883276, 7055647, 135288005, 238498066,
              229228230, 148662095, 216143425, 181639510, 101839787, 256040960, 265950570, 240677074,
              85922744, 123185272, 254450415, 97765534, 10571783, 170227406, 14542514, 40475021,
              117496916, 193371292, 250166212, 167885779, 192696288, 159404461, 130557622, 37051834,
              106640438, 183348420, 234030247, 41155851, 90597117, 173702965, 209086118, 258612781,
              189881206, 186592442, 10130658, 139182289, 241125460, 243304319, 176471684, 83853696,
              209161759, 236144340, 231358848, 230433664, 245906264, 189591954, 63350037, 54284329,
              55721255, 254509489, 47751177, 15417588, 64217206, 66148505, 229216409, 108083129,
              40553702, 118518376, 204666342, 241682233, 214551729, 108810259, 33479018, 223427563,
              226739459, 67012048, 34119889, 77337691, 246744565, 104174682, 2795054, 161827885,
              104557084, 155168409, 96142103, 118841873, 104784816, 3883583, 41086336, 134866823,
              122008382, 25569479, 211668928, 123954975, 225636920, 120936039, 197074908, 210298252,
              47994339, 13519489, 252442032, 162031725, 168407516, 132703565, 9720223, 19493867,
              184226747, 71933862, 143969713, 230702770, 69161747, 180525688, 245828202, 13250338,
              239545014, 139555205, 98878775, 9446767, 72738487, 171721518, 217644581, 249970613}))
  stage_4_butterfly_9 (
    .x_in(stage_3_per_out[18]),
    .y_in(stage_3_per_out[19]),
    .x_out(stage_4_per_in[18]),
    .y_out(stage_4_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 261793746, 116401819, 18729522, 11101448, 68136911, 71064168, 166886297,
              189762285, 21713495, 81956368, 176917280, 244883276, 7055647, 135288005, 238498066,
              229228230, 148662095, 216143425, 181639510, 101839787, 256040960, 265950570, 240677074,
              85922744, 123185272, 254450415, 97765534, 10571783, 170227406, 14542514, 40475021,
              117496916, 193371292, 250166212, 167885779, 192696288, 159404461, 130557622, 37051834,
              106640438, 183348420, 234030247, 41155851, 90597117, 173702965, 209086118, 258612781,
              189881206, 186592442, 10130658, 139182289, 241125460, 243304319, 176471684, 83853696,
              209161759, 236144340, 231358848, 230433664, 245906264, 189591954, 63350037, 54284329,
              55721255, 254509489, 47751177, 15417588, 64217206, 66148505, 229216409, 108083129,
              40553702, 118518376, 204666342, 241682233, 214551729, 108810259, 33479018, 223427563,
              226739459, 67012048, 34119889, 77337691, 246744565, 104174682, 2795054, 161827885,
              104557084, 155168409, 96142103, 118841873, 104784816, 3883583, 41086336, 134866823,
              122008382, 25569479, 211668928, 123954975, 225636920, 120936039, 197074908, 210298252,
              47994339, 13519489, 252442032, 162031725, 168407516, 132703565, 9720223, 19493867,
              184226747, 71933862, 143969713, 230702770, 69161747, 180525688, 245828202, 13250338,
              239545014, 139555205, 98878775, 9446767, 72738487, 171721518, 217644581, 249970613}))
  stage_4_butterfly_10 (
    .x_in(stage_3_per_out[20]),
    .y_in(stage_3_per_out[21]),
    .x_out(stage_4_per_in[20]),
    .y_out(stage_4_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 261793746, 116401819, 18729522, 11101448, 68136911, 71064168, 166886297,
              189762285, 21713495, 81956368, 176917280, 244883276, 7055647, 135288005, 238498066,
              229228230, 148662095, 216143425, 181639510, 101839787, 256040960, 265950570, 240677074,
              85922744, 123185272, 254450415, 97765534, 10571783, 170227406, 14542514, 40475021,
              117496916, 193371292, 250166212, 167885779, 192696288, 159404461, 130557622, 37051834,
              106640438, 183348420, 234030247, 41155851, 90597117, 173702965, 209086118, 258612781,
              189881206, 186592442, 10130658, 139182289, 241125460, 243304319, 176471684, 83853696,
              209161759, 236144340, 231358848, 230433664, 245906264, 189591954, 63350037, 54284329,
              55721255, 254509489, 47751177, 15417588, 64217206, 66148505, 229216409, 108083129,
              40553702, 118518376, 204666342, 241682233, 214551729, 108810259, 33479018, 223427563,
              226739459, 67012048, 34119889, 77337691, 246744565, 104174682, 2795054, 161827885,
              104557084, 155168409, 96142103, 118841873, 104784816, 3883583, 41086336, 134866823,
              122008382, 25569479, 211668928, 123954975, 225636920, 120936039, 197074908, 210298252,
              47994339, 13519489, 252442032, 162031725, 168407516, 132703565, 9720223, 19493867,
              184226747, 71933862, 143969713, 230702770, 69161747, 180525688, 245828202, 13250338,
              239545014, 139555205, 98878775, 9446767, 72738487, 171721518, 217644581, 249970613}))
  stage_4_butterfly_11 (
    .x_in(stage_3_per_out[22]),
    .y_in(stage_3_per_out[23]),
    .x_out(stage_4_per_in[22]),
    .y_out(stage_4_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 261793746, 116401819, 18729522, 11101448, 68136911, 71064168, 166886297,
              189762285, 21713495, 81956368, 176917280, 244883276, 7055647, 135288005, 238498066,
              229228230, 148662095, 216143425, 181639510, 101839787, 256040960, 265950570, 240677074,
              85922744, 123185272, 254450415, 97765534, 10571783, 170227406, 14542514, 40475021,
              117496916, 193371292, 250166212, 167885779, 192696288, 159404461, 130557622, 37051834,
              106640438, 183348420, 234030247, 41155851, 90597117, 173702965, 209086118, 258612781,
              189881206, 186592442, 10130658, 139182289, 241125460, 243304319, 176471684, 83853696,
              209161759, 236144340, 231358848, 230433664, 245906264, 189591954, 63350037, 54284329,
              55721255, 254509489, 47751177, 15417588, 64217206, 66148505, 229216409, 108083129,
              40553702, 118518376, 204666342, 241682233, 214551729, 108810259, 33479018, 223427563,
              226739459, 67012048, 34119889, 77337691, 246744565, 104174682, 2795054, 161827885,
              104557084, 155168409, 96142103, 118841873, 104784816, 3883583, 41086336, 134866823,
              122008382, 25569479, 211668928, 123954975, 225636920, 120936039, 197074908, 210298252,
              47994339, 13519489, 252442032, 162031725, 168407516, 132703565, 9720223, 19493867,
              184226747, 71933862, 143969713, 230702770, 69161747, 180525688, 245828202, 13250338,
              239545014, 139555205, 98878775, 9446767, 72738487, 171721518, 217644581, 249970613}))
  stage_4_butterfly_12 (
    .x_in(stage_3_per_out[24]),
    .y_in(stage_3_per_out[25]),
    .x_out(stage_4_per_in[24]),
    .y_out(stage_4_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 261793746, 116401819, 18729522, 11101448, 68136911, 71064168, 166886297,
              189762285, 21713495, 81956368, 176917280, 244883276, 7055647, 135288005, 238498066,
              229228230, 148662095, 216143425, 181639510, 101839787, 256040960, 265950570, 240677074,
              85922744, 123185272, 254450415, 97765534, 10571783, 170227406, 14542514, 40475021,
              117496916, 193371292, 250166212, 167885779, 192696288, 159404461, 130557622, 37051834,
              106640438, 183348420, 234030247, 41155851, 90597117, 173702965, 209086118, 258612781,
              189881206, 186592442, 10130658, 139182289, 241125460, 243304319, 176471684, 83853696,
              209161759, 236144340, 231358848, 230433664, 245906264, 189591954, 63350037, 54284329,
              55721255, 254509489, 47751177, 15417588, 64217206, 66148505, 229216409, 108083129,
              40553702, 118518376, 204666342, 241682233, 214551729, 108810259, 33479018, 223427563,
              226739459, 67012048, 34119889, 77337691, 246744565, 104174682, 2795054, 161827885,
              104557084, 155168409, 96142103, 118841873, 104784816, 3883583, 41086336, 134866823,
              122008382, 25569479, 211668928, 123954975, 225636920, 120936039, 197074908, 210298252,
              47994339, 13519489, 252442032, 162031725, 168407516, 132703565, 9720223, 19493867,
              184226747, 71933862, 143969713, 230702770, 69161747, 180525688, 245828202, 13250338,
              239545014, 139555205, 98878775, 9446767, 72738487, 171721518, 217644581, 249970613}))
  stage_4_butterfly_13 (
    .x_in(stage_3_per_out[26]),
    .y_in(stage_3_per_out[27]),
    .x_out(stage_4_per_in[26]),
    .y_out(stage_4_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 261793746, 116401819, 18729522, 11101448, 68136911, 71064168, 166886297,
              189762285, 21713495, 81956368, 176917280, 244883276, 7055647, 135288005, 238498066,
              229228230, 148662095, 216143425, 181639510, 101839787, 256040960, 265950570, 240677074,
              85922744, 123185272, 254450415, 97765534, 10571783, 170227406, 14542514, 40475021,
              117496916, 193371292, 250166212, 167885779, 192696288, 159404461, 130557622, 37051834,
              106640438, 183348420, 234030247, 41155851, 90597117, 173702965, 209086118, 258612781,
              189881206, 186592442, 10130658, 139182289, 241125460, 243304319, 176471684, 83853696,
              209161759, 236144340, 231358848, 230433664, 245906264, 189591954, 63350037, 54284329,
              55721255, 254509489, 47751177, 15417588, 64217206, 66148505, 229216409, 108083129,
              40553702, 118518376, 204666342, 241682233, 214551729, 108810259, 33479018, 223427563,
              226739459, 67012048, 34119889, 77337691, 246744565, 104174682, 2795054, 161827885,
              104557084, 155168409, 96142103, 118841873, 104784816, 3883583, 41086336, 134866823,
              122008382, 25569479, 211668928, 123954975, 225636920, 120936039, 197074908, 210298252,
              47994339, 13519489, 252442032, 162031725, 168407516, 132703565, 9720223, 19493867,
              184226747, 71933862, 143969713, 230702770, 69161747, 180525688, 245828202, 13250338,
              239545014, 139555205, 98878775, 9446767, 72738487, 171721518, 217644581, 249970613}))
  stage_4_butterfly_14 (
    .x_in(stage_3_per_out[28]),
    .y_in(stage_3_per_out[29]),
    .x_out(stage_4_per_in[28]),
    .y_out(stage_4_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[4]),
    .factors({80159028, 261793746, 116401819, 18729522, 11101448, 68136911, 71064168, 166886297,
              189762285, 21713495, 81956368, 176917280, 244883276, 7055647, 135288005, 238498066,
              229228230, 148662095, 216143425, 181639510, 101839787, 256040960, 265950570, 240677074,
              85922744, 123185272, 254450415, 97765534, 10571783, 170227406, 14542514, 40475021,
              117496916, 193371292, 250166212, 167885779, 192696288, 159404461, 130557622, 37051834,
              106640438, 183348420, 234030247, 41155851, 90597117, 173702965, 209086118, 258612781,
              189881206, 186592442, 10130658, 139182289, 241125460, 243304319, 176471684, 83853696,
              209161759, 236144340, 231358848, 230433664, 245906264, 189591954, 63350037, 54284329,
              55721255, 254509489, 47751177, 15417588, 64217206, 66148505, 229216409, 108083129,
              40553702, 118518376, 204666342, 241682233, 214551729, 108810259, 33479018, 223427563,
              226739459, 67012048, 34119889, 77337691, 246744565, 104174682, 2795054, 161827885,
              104557084, 155168409, 96142103, 118841873, 104784816, 3883583, 41086336, 134866823,
              122008382, 25569479, 211668928, 123954975, 225636920, 120936039, 197074908, 210298252,
              47994339, 13519489, 252442032, 162031725, 168407516, 132703565, 9720223, 19493867,
              184226747, 71933862, 143969713, 230702770, 69161747, 180525688, 245828202, 13250338,
              239545014, 139555205, 98878775, 9446767, 72738487, 171721518, 217644581, 249970613}))
  stage_4_butterfly_15 (
    .x_in(stage_3_per_out[30]),
    .y_in(stage_3_per_out[31]),
    .x_out(stage_4_per_in[30]),
    .y_out(stage_4_per_in[31]),
    .clk(clk),
    .rst(rst)
  );





  // TODO(Yang): stage 4 -> stage 5 permutation
  // FIXME: ignore butterfly units for now.
  stage_4_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_4_5_per (
    .inData_0(stage_4_per_in[0]),
    .inData_1(stage_4_per_in[1]),
    .inData_2(stage_4_per_in[2]),
    .inData_3(stage_4_per_in[3]),
    .inData_4(stage_4_per_in[4]),
    .inData_5(stage_4_per_in[5]),
    .inData_6(stage_4_per_in[6]),
    .inData_7(stage_4_per_in[7]),
    .inData_8(stage_4_per_in[8]),
    .inData_9(stage_4_per_in[9]),
    .inData_10(stage_4_per_in[10]),
    .inData_11(stage_4_per_in[11]),
    .inData_12(stage_4_per_in[12]),
    .inData_13(stage_4_per_in[13]),
    .inData_14(stage_4_per_in[14]),
    .inData_15(stage_4_per_in[15]),
    .inData_16(stage_4_per_in[16]),
    .inData_17(stage_4_per_in[17]),
    .inData_18(stage_4_per_in[18]),
    .inData_19(stage_4_per_in[19]),
    .inData_20(stage_4_per_in[20]),
    .inData_21(stage_4_per_in[21]),
    .inData_22(stage_4_per_in[22]),
    .inData_23(stage_4_per_in[23]),
    .inData_24(stage_4_per_in[24]),
    .inData_25(stage_4_per_in[25]),
    .inData_26(stage_4_per_in[26]),
    .inData_27(stage_4_per_in[27]),
    .inData_28(stage_4_per_in[28]),
    .inData_29(stage_4_per_in[29]),
    .inData_30(stage_4_per_in[30]),
    .inData_31(stage_4_per_in[31]),
    .outData_0(stage_4_per_out[0]),
    .outData_1(stage_4_per_out[1]),
    .outData_2(stage_4_per_out[2]),
    .outData_3(stage_4_per_out[3]),
    .outData_4(stage_4_per_out[4]),
    .outData_5(stage_4_per_out[5]),
    .outData_6(stage_4_per_out[6]),
    .outData_7(stage_4_per_out[7]),
    .outData_8(stage_4_per_out[8]),
    .outData_9(stage_4_per_out[9]),
    .outData_10(stage_4_per_out[10]),
    .outData_11(stage_4_per_out[11]),
    .outData_12(stage_4_per_out[12]),
    .outData_13(stage_4_per_out[13]),
    .outData_14(stage_4_per_out[14]),
    .outData_15(stage_4_per_out[15]),
    .outData_16(stage_4_per_out[16]),
    .outData_17(stage_4_per_out[17]),
    .outData_18(stage_4_per_out[18]),
    .outData_19(stage_4_per_out[19]),
    .outData_20(stage_4_per_out[20]),
    .outData_21(stage_4_per_out[21]),
    .outData_22(stage_4_per_out[22]),
    .outData_23(stage_4_per_out[23]),
    .outData_24(stage_4_per_out[24]),
    .outData_25(stage_4_per_out[25]),
    .outData_26(stage_4_per_out[26]),
    .outData_27(stage_4_per_out[27]),
    .outData_28(stage_4_per_out[28]),
    .outData_29(stage_4_per_out[29]),
    .outData_30(stage_4_per_out[30]),
    .outData_31(stage_4_per_out[31]),
    .in_start(in_start[4]),
    .out_start(out_start[4]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 5 32 butterfly units
  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 124918999, 185598009, 185598009, 239095400, 239095400, 39593842, 39593842,
              169276669, 169276669, 141548072, 141548072, 197386970, 197386970, 119224607, 119224607,
              159115155, 159115155, 208403048, 208403048, 102065274, 102065274, 111284191, 111284191,
              157028693, 157028693, 30748955, 30748955, 210568560, 210568560, 91114882, 91114882,
              74680748, 74680748, 162373432, 162373432, 155896930, 155896930, 145384235, 145384235,
              100099056, 100099056, 71471012, 71471012, 136571165, 136571165, 33165861, 33165861,
              149429971, 149429971, 206324144, 206324144, 175609590, 175609590, 152865265, 152865265,
              201062854, 201062854, 138074788, 138074788, 191727270, 191727270, 41084242, 41084242,
              227611463, 227611463, 196909902, 196909902, 49823188, 49823188, 78852289, 78852289,
              202366126, 202366126, 146694818, 146694818, 120670867, 120670867, 86517113, 86517113,
              256674305, 256674305, 114407843, 114407843, 233560477, 233560477, 78462606, 78462606,
              92577793, 92577793, 70582130, 70582130, 172642311, 172642311, 215696667, 215696667,
              251290023, 251290023, 193045667, 193045667, 202257393, 202257393, 242795574, 242795574,
              240684902, 240684902, 47317233, 47317233, 263678998, 263678998, 152412548, 152412548,
              200054106, 200054106, 76707105, 76707105, 140204941, 140204941, 170752771, 170752771,
              109553202, 109553202, 179817683, 179817683, 262046585, 262046585, 165226744, 165226744}))
  stage_5_butterfly_0 (
    .x_in(stage_4_per_out[0]),
    .y_in(stage_4_per_out[1]),
    .x_out(stage_5_per_in[0]),
    .y_out(stage_5_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 124918999, 185598009, 185598009, 239095400, 239095400, 39593842, 39593842,
              169276669, 169276669, 141548072, 141548072, 197386970, 197386970, 119224607, 119224607,
              159115155, 159115155, 208403048, 208403048, 102065274, 102065274, 111284191, 111284191,
              157028693, 157028693, 30748955, 30748955, 210568560, 210568560, 91114882, 91114882,
              74680748, 74680748, 162373432, 162373432, 155896930, 155896930, 145384235, 145384235,
              100099056, 100099056, 71471012, 71471012, 136571165, 136571165, 33165861, 33165861,
              149429971, 149429971, 206324144, 206324144, 175609590, 175609590, 152865265, 152865265,
              201062854, 201062854, 138074788, 138074788, 191727270, 191727270, 41084242, 41084242,
              227611463, 227611463, 196909902, 196909902, 49823188, 49823188, 78852289, 78852289,
              202366126, 202366126, 146694818, 146694818, 120670867, 120670867, 86517113, 86517113,
              256674305, 256674305, 114407843, 114407843, 233560477, 233560477, 78462606, 78462606,
              92577793, 92577793, 70582130, 70582130, 172642311, 172642311, 215696667, 215696667,
              251290023, 251290023, 193045667, 193045667, 202257393, 202257393, 242795574, 242795574,
              240684902, 240684902, 47317233, 47317233, 263678998, 263678998, 152412548, 152412548,
              200054106, 200054106, 76707105, 76707105, 140204941, 140204941, 170752771, 170752771,
              109553202, 109553202, 179817683, 179817683, 262046585, 262046585, 165226744, 165226744}))
  stage_5_butterfly_1 (
    .x_in(stage_4_per_out[2]),
    .y_in(stage_4_per_out[3]),
    .x_out(stage_5_per_in[2]),
    .y_out(stage_5_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 124918999, 185598009, 185598009, 239095400, 239095400, 39593842, 39593842,
              169276669, 169276669, 141548072, 141548072, 197386970, 197386970, 119224607, 119224607,
              159115155, 159115155, 208403048, 208403048, 102065274, 102065274, 111284191, 111284191,
              157028693, 157028693, 30748955, 30748955, 210568560, 210568560, 91114882, 91114882,
              74680748, 74680748, 162373432, 162373432, 155896930, 155896930, 145384235, 145384235,
              100099056, 100099056, 71471012, 71471012, 136571165, 136571165, 33165861, 33165861,
              149429971, 149429971, 206324144, 206324144, 175609590, 175609590, 152865265, 152865265,
              201062854, 201062854, 138074788, 138074788, 191727270, 191727270, 41084242, 41084242,
              227611463, 227611463, 196909902, 196909902, 49823188, 49823188, 78852289, 78852289,
              202366126, 202366126, 146694818, 146694818, 120670867, 120670867, 86517113, 86517113,
              256674305, 256674305, 114407843, 114407843, 233560477, 233560477, 78462606, 78462606,
              92577793, 92577793, 70582130, 70582130, 172642311, 172642311, 215696667, 215696667,
              251290023, 251290023, 193045667, 193045667, 202257393, 202257393, 242795574, 242795574,
              240684902, 240684902, 47317233, 47317233, 263678998, 263678998, 152412548, 152412548,
              200054106, 200054106, 76707105, 76707105, 140204941, 140204941, 170752771, 170752771,
              109553202, 109553202, 179817683, 179817683, 262046585, 262046585, 165226744, 165226744}))
  stage_5_butterfly_2 (
    .x_in(stage_4_per_out[4]),
    .y_in(stage_4_per_out[5]),
    .x_out(stage_5_per_in[4]),
    .y_out(stage_5_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 124918999, 185598009, 185598009, 239095400, 239095400, 39593842, 39593842,
              169276669, 169276669, 141548072, 141548072, 197386970, 197386970, 119224607, 119224607,
              159115155, 159115155, 208403048, 208403048, 102065274, 102065274, 111284191, 111284191,
              157028693, 157028693, 30748955, 30748955, 210568560, 210568560, 91114882, 91114882,
              74680748, 74680748, 162373432, 162373432, 155896930, 155896930, 145384235, 145384235,
              100099056, 100099056, 71471012, 71471012, 136571165, 136571165, 33165861, 33165861,
              149429971, 149429971, 206324144, 206324144, 175609590, 175609590, 152865265, 152865265,
              201062854, 201062854, 138074788, 138074788, 191727270, 191727270, 41084242, 41084242,
              227611463, 227611463, 196909902, 196909902, 49823188, 49823188, 78852289, 78852289,
              202366126, 202366126, 146694818, 146694818, 120670867, 120670867, 86517113, 86517113,
              256674305, 256674305, 114407843, 114407843, 233560477, 233560477, 78462606, 78462606,
              92577793, 92577793, 70582130, 70582130, 172642311, 172642311, 215696667, 215696667,
              251290023, 251290023, 193045667, 193045667, 202257393, 202257393, 242795574, 242795574,
              240684902, 240684902, 47317233, 47317233, 263678998, 263678998, 152412548, 152412548,
              200054106, 200054106, 76707105, 76707105, 140204941, 140204941, 170752771, 170752771,
              109553202, 109553202, 179817683, 179817683, 262046585, 262046585, 165226744, 165226744}))
  stage_5_butterfly_3 (
    .x_in(stage_4_per_out[6]),
    .y_in(stage_4_per_out[7]),
    .x_out(stage_5_per_in[6]),
    .y_out(stage_5_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 124918999, 185598009, 185598009, 239095400, 239095400, 39593842, 39593842,
              169276669, 169276669, 141548072, 141548072, 197386970, 197386970, 119224607, 119224607,
              159115155, 159115155, 208403048, 208403048, 102065274, 102065274, 111284191, 111284191,
              157028693, 157028693, 30748955, 30748955, 210568560, 210568560, 91114882, 91114882,
              74680748, 74680748, 162373432, 162373432, 155896930, 155896930, 145384235, 145384235,
              100099056, 100099056, 71471012, 71471012, 136571165, 136571165, 33165861, 33165861,
              149429971, 149429971, 206324144, 206324144, 175609590, 175609590, 152865265, 152865265,
              201062854, 201062854, 138074788, 138074788, 191727270, 191727270, 41084242, 41084242,
              227611463, 227611463, 196909902, 196909902, 49823188, 49823188, 78852289, 78852289,
              202366126, 202366126, 146694818, 146694818, 120670867, 120670867, 86517113, 86517113,
              256674305, 256674305, 114407843, 114407843, 233560477, 233560477, 78462606, 78462606,
              92577793, 92577793, 70582130, 70582130, 172642311, 172642311, 215696667, 215696667,
              251290023, 251290023, 193045667, 193045667, 202257393, 202257393, 242795574, 242795574,
              240684902, 240684902, 47317233, 47317233, 263678998, 263678998, 152412548, 152412548,
              200054106, 200054106, 76707105, 76707105, 140204941, 140204941, 170752771, 170752771,
              109553202, 109553202, 179817683, 179817683, 262046585, 262046585, 165226744, 165226744}))
  stage_5_butterfly_4 (
    .x_in(stage_4_per_out[8]),
    .y_in(stage_4_per_out[9]),
    .x_out(stage_5_per_in[8]),
    .y_out(stage_5_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 124918999, 185598009, 185598009, 239095400, 239095400, 39593842, 39593842,
              169276669, 169276669, 141548072, 141548072, 197386970, 197386970, 119224607, 119224607,
              159115155, 159115155, 208403048, 208403048, 102065274, 102065274, 111284191, 111284191,
              157028693, 157028693, 30748955, 30748955, 210568560, 210568560, 91114882, 91114882,
              74680748, 74680748, 162373432, 162373432, 155896930, 155896930, 145384235, 145384235,
              100099056, 100099056, 71471012, 71471012, 136571165, 136571165, 33165861, 33165861,
              149429971, 149429971, 206324144, 206324144, 175609590, 175609590, 152865265, 152865265,
              201062854, 201062854, 138074788, 138074788, 191727270, 191727270, 41084242, 41084242,
              227611463, 227611463, 196909902, 196909902, 49823188, 49823188, 78852289, 78852289,
              202366126, 202366126, 146694818, 146694818, 120670867, 120670867, 86517113, 86517113,
              256674305, 256674305, 114407843, 114407843, 233560477, 233560477, 78462606, 78462606,
              92577793, 92577793, 70582130, 70582130, 172642311, 172642311, 215696667, 215696667,
              251290023, 251290023, 193045667, 193045667, 202257393, 202257393, 242795574, 242795574,
              240684902, 240684902, 47317233, 47317233, 263678998, 263678998, 152412548, 152412548,
              200054106, 200054106, 76707105, 76707105, 140204941, 140204941, 170752771, 170752771,
              109553202, 109553202, 179817683, 179817683, 262046585, 262046585, 165226744, 165226744}))
  stage_5_butterfly_5 (
    .x_in(stage_4_per_out[10]),
    .y_in(stage_4_per_out[11]),
    .x_out(stage_5_per_in[10]),
    .y_out(stage_5_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 124918999, 185598009, 185598009, 239095400, 239095400, 39593842, 39593842,
              169276669, 169276669, 141548072, 141548072, 197386970, 197386970, 119224607, 119224607,
              159115155, 159115155, 208403048, 208403048, 102065274, 102065274, 111284191, 111284191,
              157028693, 157028693, 30748955, 30748955, 210568560, 210568560, 91114882, 91114882,
              74680748, 74680748, 162373432, 162373432, 155896930, 155896930, 145384235, 145384235,
              100099056, 100099056, 71471012, 71471012, 136571165, 136571165, 33165861, 33165861,
              149429971, 149429971, 206324144, 206324144, 175609590, 175609590, 152865265, 152865265,
              201062854, 201062854, 138074788, 138074788, 191727270, 191727270, 41084242, 41084242,
              227611463, 227611463, 196909902, 196909902, 49823188, 49823188, 78852289, 78852289,
              202366126, 202366126, 146694818, 146694818, 120670867, 120670867, 86517113, 86517113,
              256674305, 256674305, 114407843, 114407843, 233560477, 233560477, 78462606, 78462606,
              92577793, 92577793, 70582130, 70582130, 172642311, 172642311, 215696667, 215696667,
              251290023, 251290023, 193045667, 193045667, 202257393, 202257393, 242795574, 242795574,
              240684902, 240684902, 47317233, 47317233, 263678998, 263678998, 152412548, 152412548,
              200054106, 200054106, 76707105, 76707105, 140204941, 140204941, 170752771, 170752771,
              109553202, 109553202, 179817683, 179817683, 262046585, 262046585, 165226744, 165226744}))
  stage_5_butterfly_6 (
    .x_in(stage_4_per_out[12]),
    .y_in(stage_4_per_out[13]),
    .x_out(stage_5_per_in[12]),
    .y_out(stage_5_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 124918999, 185598009, 185598009, 239095400, 239095400, 39593842, 39593842,
              169276669, 169276669, 141548072, 141548072, 197386970, 197386970, 119224607, 119224607,
              159115155, 159115155, 208403048, 208403048, 102065274, 102065274, 111284191, 111284191,
              157028693, 157028693, 30748955, 30748955, 210568560, 210568560, 91114882, 91114882,
              74680748, 74680748, 162373432, 162373432, 155896930, 155896930, 145384235, 145384235,
              100099056, 100099056, 71471012, 71471012, 136571165, 136571165, 33165861, 33165861,
              149429971, 149429971, 206324144, 206324144, 175609590, 175609590, 152865265, 152865265,
              201062854, 201062854, 138074788, 138074788, 191727270, 191727270, 41084242, 41084242,
              227611463, 227611463, 196909902, 196909902, 49823188, 49823188, 78852289, 78852289,
              202366126, 202366126, 146694818, 146694818, 120670867, 120670867, 86517113, 86517113,
              256674305, 256674305, 114407843, 114407843, 233560477, 233560477, 78462606, 78462606,
              92577793, 92577793, 70582130, 70582130, 172642311, 172642311, 215696667, 215696667,
              251290023, 251290023, 193045667, 193045667, 202257393, 202257393, 242795574, 242795574,
              240684902, 240684902, 47317233, 47317233, 263678998, 263678998, 152412548, 152412548,
              200054106, 200054106, 76707105, 76707105, 140204941, 140204941, 170752771, 170752771,
              109553202, 109553202, 179817683, 179817683, 262046585, 262046585, 165226744, 165226744}))
  stage_5_butterfly_7 (
    .x_in(stage_4_per_out[14]),
    .y_in(stage_4_per_out[15]),
    .x_out(stage_5_per_in[14]),
    .y_out(stage_5_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 124918999, 185598009, 185598009, 239095400, 239095400, 39593842, 39593842,
              169276669, 169276669, 141548072, 141548072, 197386970, 197386970, 119224607, 119224607,
              159115155, 159115155, 208403048, 208403048, 102065274, 102065274, 111284191, 111284191,
              157028693, 157028693, 30748955, 30748955, 210568560, 210568560, 91114882, 91114882,
              74680748, 74680748, 162373432, 162373432, 155896930, 155896930, 145384235, 145384235,
              100099056, 100099056, 71471012, 71471012, 136571165, 136571165, 33165861, 33165861,
              149429971, 149429971, 206324144, 206324144, 175609590, 175609590, 152865265, 152865265,
              201062854, 201062854, 138074788, 138074788, 191727270, 191727270, 41084242, 41084242,
              227611463, 227611463, 196909902, 196909902, 49823188, 49823188, 78852289, 78852289,
              202366126, 202366126, 146694818, 146694818, 120670867, 120670867, 86517113, 86517113,
              256674305, 256674305, 114407843, 114407843, 233560477, 233560477, 78462606, 78462606,
              92577793, 92577793, 70582130, 70582130, 172642311, 172642311, 215696667, 215696667,
              251290023, 251290023, 193045667, 193045667, 202257393, 202257393, 242795574, 242795574,
              240684902, 240684902, 47317233, 47317233, 263678998, 263678998, 152412548, 152412548,
              200054106, 200054106, 76707105, 76707105, 140204941, 140204941, 170752771, 170752771,
              109553202, 109553202, 179817683, 179817683, 262046585, 262046585, 165226744, 165226744}))
  stage_5_butterfly_8 (
    .x_in(stage_4_per_out[16]),
    .y_in(stage_4_per_out[17]),
    .x_out(stage_5_per_in[16]),
    .y_out(stage_5_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 124918999, 185598009, 185598009, 239095400, 239095400, 39593842, 39593842,
              169276669, 169276669, 141548072, 141548072, 197386970, 197386970, 119224607, 119224607,
              159115155, 159115155, 208403048, 208403048, 102065274, 102065274, 111284191, 111284191,
              157028693, 157028693, 30748955, 30748955, 210568560, 210568560, 91114882, 91114882,
              74680748, 74680748, 162373432, 162373432, 155896930, 155896930, 145384235, 145384235,
              100099056, 100099056, 71471012, 71471012, 136571165, 136571165, 33165861, 33165861,
              149429971, 149429971, 206324144, 206324144, 175609590, 175609590, 152865265, 152865265,
              201062854, 201062854, 138074788, 138074788, 191727270, 191727270, 41084242, 41084242,
              227611463, 227611463, 196909902, 196909902, 49823188, 49823188, 78852289, 78852289,
              202366126, 202366126, 146694818, 146694818, 120670867, 120670867, 86517113, 86517113,
              256674305, 256674305, 114407843, 114407843, 233560477, 233560477, 78462606, 78462606,
              92577793, 92577793, 70582130, 70582130, 172642311, 172642311, 215696667, 215696667,
              251290023, 251290023, 193045667, 193045667, 202257393, 202257393, 242795574, 242795574,
              240684902, 240684902, 47317233, 47317233, 263678998, 263678998, 152412548, 152412548,
              200054106, 200054106, 76707105, 76707105, 140204941, 140204941, 170752771, 170752771,
              109553202, 109553202, 179817683, 179817683, 262046585, 262046585, 165226744, 165226744}))
  stage_5_butterfly_9 (
    .x_in(stage_4_per_out[18]),
    .y_in(stage_4_per_out[19]),
    .x_out(stage_5_per_in[18]),
    .y_out(stage_5_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 124918999, 185598009, 185598009, 239095400, 239095400, 39593842, 39593842,
              169276669, 169276669, 141548072, 141548072, 197386970, 197386970, 119224607, 119224607,
              159115155, 159115155, 208403048, 208403048, 102065274, 102065274, 111284191, 111284191,
              157028693, 157028693, 30748955, 30748955, 210568560, 210568560, 91114882, 91114882,
              74680748, 74680748, 162373432, 162373432, 155896930, 155896930, 145384235, 145384235,
              100099056, 100099056, 71471012, 71471012, 136571165, 136571165, 33165861, 33165861,
              149429971, 149429971, 206324144, 206324144, 175609590, 175609590, 152865265, 152865265,
              201062854, 201062854, 138074788, 138074788, 191727270, 191727270, 41084242, 41084242,
              227611463, 227611463, 196909902, 196909902, 49823188, 49823188, 78852289, 78852289,
              202366126, 202366126, 146694818, 146694818, 120670867, 120670867, 86517113, 86517113,
              256674305, 256674305, 114407843, 114407843, 233560477, 233560477, 78462606, 78462606,
              92577793, 92577793, 70582130, 70582130, 172642311, 172642311, 215696667, 215696667,
              251290023, 251290023, 193045667, 193045667, 202257393, 202257393, 242795574, 242795574,
              240684902, 240684902, 47317233, 47317233, 263678998, 263678998, 152412548, 152412548,
              200054106, 200054106, 76707105, 76707105, 140204941, 140204941, 170752771, 170752771,
              109553202, 109553202, 179817683, 179817683, 262046585, 262046585, 165226744, 165226744}))
  stage_5_butterfly_10 (
    .x_in(stage_4_per_out[20]),
    .y_in(stage_4_per_out[21]),
    .x_out(stage_5_per_in[20]),
    .y_out(stage_5_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 124918999, 185598009, 185598009, 239095400, 239095400, 39593842, 39593842,
              169276669, 169276669, 141548072, 141548072, 197386970, 197386970, 119224607, 119224607,
              159115155, 159115155, 208403048, 208403048, 102065274, 102065274, 111284191, 111284191,
              157028693, 157028693, 30748955, 30748955, 210568560, 210568560, 91114882, 91114882,
              74680748, 74680748, 162373432, 162373432, 155896930, 155896930, 145384235, 145384235,
              100099056, 100099056, 71471012, 71471012, 136571165, 136571165, 33165861, 33165861,
              149429971, 149429971, 206324144, 206324144, 175609590, 175609590, 152865265, 152865265,
              201062854, 201062854, 138074788, 138074788, 191727270, 191727270, 41084242, 41084242,
              227611463, 227611463, 196909902, 196909902, 49823188, 49823188, 78852289, 78852289,
              202366126, 202366126, 146694818, 146694818, 120670867, 120670867, 86517113, 86517113,
              256674305, 256674305, 114407843, 114407843, 233560477, 233560477, 78462606, 78462606,
              92577793, 92577793, 70582130, 70582130, 172642311, 172642311, 215696667, 215696667,
              251290023, 251290023, 193045667, 193045667, 202257393, 202257393, 242795574, 242795574,
              240684902, 240684902, 47317233, 47317233, 263678998, 263678998, 152412548, 152412548,
              200054106, 200054106, 76707105, 76707105, 140204941, 140204941, 170752771, 170752771,
              109553202, 109553202, 179817683, 179817683, 262046585, 262046585, 165226744, 165226744}))
  stage_5_butterfly_11 (
    .x_in(stage_4_per_out[22]),
    .y_in(stage_4_per_out[23]),
    .x_out(stage_5_per_in[22]),
    .y_out(stage_5_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 124918999, 185598009, 185598009, 239095400, 239095400, 39593842, 39593842,
              169276669, 169276669, 141548072, 141548072, 197386970, 197386970, 119224607, 119224607,
              159115155, 159115155, 208403048, 208403048, 102065274, 102065274, 111284191, 111284191,
              157028693, 157028693, 30748955, 30748955, 210568560, 210568560, 91114882, 91114882,
              74680748, 74680748, 162373432, 162373432, 155896930, 155896930, 145384235, 145384235,
              100099056, 100099056, 71471012, 71471012, 136571165, 136571165, 33165861, 33165861,
              149429971, 149429971, 206324144, 206324144, 175609590, 175609590, 152865265, 152865265,
              201062854, 201062854, 138074788, 138074788, 191727270, 191727270, 41084242, 41084242,
              227611463, 227611463, 196909902, 196909902, 49823188, 49823188, 78852289, 78852289,
              202366126, 202366126, 146694818, 146694818, 120670867, 120670867, 86517113, 86517113,
              256674305, 256674305, 114407843, 114407843, 233560477, 233560477, 78462606, 78462606,
              92577793, 92577793, 70582130, 70582130, 172642311, 172642311, 215696667, 215696667,
              251290023, 251290023, 193045667, 193045667, 202257393, 202257393, 242795574, 242795574,
              240684902, 240684902, 47317233, 47317233, 263678998, 263678998, 152412548, 152412548,
              200054106, 200054106, 76707105, 76707105, 140204941, 140204941, 170752771, 170752771,
              109553202, 109553202, 179817683, 179817683, 262046585, 262046585, 165226744, 165226744}))
  stage_5_butterfly_12 (
    .x_in(stage_4_per_out[24]),
    .y_in(stage_4_per_out[25]),
    .x_out(stage_5_per_in[24]),
    .y_out(stage_5_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 124918999, 185598009, 185598009, 239095400, 239095400, 39593842, 39593842,
              169276669, 169276669, 141548072, 141548072, 197386970, 197386970, 119224607, 119224607,
              159115155, 159115155, 208403048, 208403048, 102065274, 102065274, 111284191, 111284191,
              157028693, 157028693, 30748955, 30748955, 210568560, 210568560, 91114882, 91114882,
              74680748, 74680748, 162373432, 162373432, 155896930, 155896930, 145384235, 145384235,
              100099056, 100099056, 71471012, 71471012, 136571165, 136571165, 33165861, 33165861,
              149429971, 149429971, 206324144, 206324144, 175609590, 175609590, 152865265, 152865265,
              201062854, 201062854, 138074788, 138074788, 191727270, 191727270, 41084242, 41084242,
              227611463, 227611463, 196909902, 196909902, 49823188, 49823188, 78852289, 78852289,
              202366126, 202366126, 146694818, 146694818, 120670867, 120670867, 86517113, 86517113,
              256674305, 256674305, 114407843, 114407843, 233560477, 233560477, 78462606, 78462606,
              92577793, 92577793, 70582130, 70582130, 172642311, 172642311, 215696667, 215696667,
              251290023, 251290023, 193045667, 193045667, 202257393, 202257393, 242795574, 242795574,
              240684902, 240684902, 47317233, 47317233, 263678998, 263678998, 152412548, 152412548,
              200054106, 200054106, 76707105, 76707105, 140204941, 140204941, 170752771, 170752771,
              109553202, 109553202, 179817683, 179817683, 262046585, 262046585, 165226744, 165226744}))
  stage_5_butterfly_13 (
    .x_in(stage_4_per_out[26]),
    .y_in(stage_4_per_out[27]),
    .x_out(stage_5_per_in[26]),
    .y_out(stage_5_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 124918999, 185598009, 185598009, 239095400, 239095400, 39593842, 39593842,
              169276669, 169276669, 141548072, 141548072, 197386970, 197386970, 119224607, 119224607,
              159115155, 159115155, 208403048, 208403048, 102065274, 102065274, 111284191, 111284191,
              157028693, 157028693, 30748955, 30748955, 210568560, 210568560, 91114882, 91114882,
              74680748, 74680748, 162373432, 162373432, 155896930, 155896930, 145384235, 145384235,
              100099056, 100099056, 71471012, 71471012, 136571165, 136571165, 33165861, 33165861,
              149429971, 149429971, 206324144, 206324144, 175609590, 175609590, 152865265, 152865265,
              201062854, 201062854, 138074788, 138074788, 191727270, 191727270, 41084242, 41084242,
              227611463, 227611463, 196909902, 196909902, 49823188, 49823188, 78852289, 78852289,
              202366126, 202366126, 146694818, 146694818, 120670867, 120670867, 86517113, 86517113,
              256674305, 256674305, 114407843, 114407843, 233560477, 233560477, 78462606, 78462606,
              92577793, 92577793, 70582130, 70582130, 172642311, 172642311, 215696667, 215696667,
              251290023, 251290023, 193045667, 193045667, 202257393, 202257393, 242795574, 242795574,
              240684902, 240684902, 47317233, 47317233, 263678998, 263678998, 152412548, 152412548,
              200054106, 200054106, 76707105, 76707105, 140204941, 140204941, 170752771, 170752771,
              109553202, 109553202, 179817683, 179817683, 262046585, 262046585, 165226744, 165226744}))
  stage_5_butterfly_14 (
    .x_in(stage_4_per_out[28]),
    .y_in(stage_4_per_out[29]),
    .x_out(stage_5_per_in[28]),
    .y_out(stage_5_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[5]),
    .factors({124918999, 124918999, 185598009, 185598009, 239095400, 239095400, 39593842, 39593842,
              169276669, 169276669, 141548072, 141548072, 197386970, 197386970, 119224607, 119224607,
              159115155, 159115155, 208403048, 208403048, 102065274, 102065274, 111284191, 111284191,
              157028693, 157028693, 30748955, 30748955, 210568560, 210568560, 91114882, 91114882,
              74680748, 74680748, 162373432, 162373432, 155896930, 155896930, 145384235, 145384235,
              100099056, 100099056, 71471012, 71471012, 136571165, 136571165, 33165861, 33165861,
              149429971, 149429971, 206324144, 206324144, 175609590, 175609590, 152865265, 152865265,
              201062854, 201062854, 138074788, 138074788, 191727270, 191727270, 41084242, 41084242,
              227611463, 227611463, 196909902, 196909902, 49823188, 49823188, 78852289, 78852289,
              202366126, 202366126, 146694818, 146694818, 120670867, 120670867, 86517113, 86517113,
              256674305, 256674305, 114407843, 114407843, 233560477, 233560477, 78462606, 78462606,
              92577793, 92577793, 70582130, 70582130, 172642311, 172642311, 215696667, 215696667,
              251290023, 251290023, 193045667, 193045667, 202257393, 202257393, 242795574, 242795574,
              240684902, 240684902, 47317233, 47317233, 263678998, 263678998, 152412548, 152412548,
              200054106, 200054106, 76707105, 76707105, 140204941, 140204941, 170752771, 170752771,
              109553202, 109553202, 179817683, 179817683, 262046585, 262046585, 165226744, 165226744}))
  stage_5_butterfly_15 (
    .x_in(stage_4_per_out[30]),
    .y_in(stage_4_per_out[31]),
    .x_out(stage_5_per_in[30]),
    .y_out(stage_5_per_in[31]),
    .clk(clk),
    .rst(rst)
  );






  // TODO(Yang): stage 5 -> stage 6 permutation
  // FIXME: ignore butterfly units for now.
  stage_5_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_5_6_per (
    .inData_0(stage_5_per_in[0]),
    .inData_1(stage_5_per_in[1]),
    .inData_2(stage_5_per_in[2]),
    .inData_3(stage_5_per_in[3]),
    .inData_4(stage_5_per_in[4]),
    .inData_5(stage_5_per_in[5]),
    .inData_6(stage_5_per_in[6]),
    .inData_7(stage_5_per_in[7]),
    .inData_8(stage_5_per_in[8]),
    .inData_9(stage_5_per_in[9]),
    .inData_10(stage_5_per_in[10]),
    .inData_11(stage_5_per_in[11]),
    .inData_12(stage_5_per_in[12]),
    .inData_13(stage_5_per_in[13]),
    .inData_14(stage_5_per_in[14]),
    .inData_15(stage_5_per_in[15]),
    .inData_16(stage_5_per_in[16]),
    .inData_17(stage_5_per_in[17]),
    .inData_18(stage_5_per_in[18]),
    .inData_19(stage_5_per_in[19]),
    .inData_20(stage_5_per_in[20]),
    .inData_21(stage_5_per_in[21]),
    .inData_22(stage_5_per_in[22]),
    .inData_23(stage_5_per_in[23]),
    .inData_24(stage_5_per_in[24]),
    .inData_25(stage_5_per_in[25]),
    .inData_26(stage_5_per_in[26]),
    .inData_27(stage_5_per_in[27]),
    .inData_28(stage_5_per_in[28]),
    .inData_29(stage_5_per_in[29]),
    .inData_30(stage_5_per_in[30]),
    .inData_31(stage_5_per_in[31]),
    .outData_0(stage_5_per_out[0]),
    .outData_1(stage_5_per_out[1]),
    .outData_2(stage_5_per_out[2]),
    .outData_3(stage_5_per_out[3]),
    .outData_4(stage_5_per_out[4]),
    .outData_5(stage_5_per_out[5]),
    .outData_6(stage_5_per_out[6]),
    .outData_7(stage_5_per_out[7]),
    .outData_8(stage_5_per_out[8]),
    .outData_9(stage_5_per_out[9]),
    .outData_10(stage_5_per_out[10]),
    .outData_11(stage_5_per_out[11]),
    .outData_12(stage_5_per_out[12]),
    .outData_13(stage_5_per_out[13]),
    .outData_14(stage_5_per_out[14]),
    .outData_15(stage_5_per_out[15]),
    .outData_16(stage_5_per_out[16]),
    .outData_17(stage_5_per_out[17]),
    .outData_18(stage_5_per_out[18]),
    .outData_19(stage_5_per_out[19]),
    .outData_20(stage_5_per_out[20]),
    .outData_21(stage_5_per_out[21]),
    .outData_22(stage_5_per_out[22]),
    .outData_23(stage_5_per_out[23]),
    .outData_24(stage_5_per_out[24]),
    .outData_25(stage_5_per_out[25]),
    .outData_26(stage_5_per_out[26]),
    .outData_27(stage_5_per_out[27]),
    .outData_28(stage_5_per_out[28]),
    .outData_29(stage_5_per_out[29]),
    .outData_30(stage_5_per_out[30]),
    .outData_31(stage_5_per_out[31]),
    .in_start(in_start[5]),
    .out_start(out_start[5]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 6 32 butterfly units
  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 265190919, 265190919, 102773617, 102773617, 102773617, 102773617,
              210831626, 210831626, 210831626, 210831626, 84893967, 84893967, 84893967, 84893967,
              119480423, 119480423, 119480423, 119480423, 102579498, 102579498, 102579498, 102579498,
              129001811, 129001811, 129001811, 129001811, 72061017, 72061017, 72061017, 72061017,
              72052889, 72052889, 72052889, 72052889, 73825164, 73825164, 73825164, 73825164,
              18533839, 18533839, 18533839, 18533839, 168579404, 168579404, 168579404, 168579404,
              47877183, 47877183, 47877183, 47877183, 184798272, 184798272, 184798272, 184798272,
              5258704, 5258704, 5258704, 5258704, 92744225, 92744225, 92744225, 92744225,
              221840088, 221840088, 221840088, 221840088, 216372172, 216372172, 216372172, 216372172,
              231414272, 231414272, 231414272, 231414272, 94135184, 94135184, 94135184, 94135184,
              89995519, 89995519, 89995519, 89995519, 220656190, 220656190, 220656190, 220656190,
              183300662, 183300662, 183300662, 183300662, 160020761, 160020761, 160020761, 160020761,
              249274747, 249274747, 249274747, 249274747, 62061822, 62061822, 62061822, 62061822,
              76573097, 76573097, 76573097, 76573097, 35289455, 35289455, 35289455, 35289455,
              234642902, 234642902, 234642902, 234642902, 229105823, 229105823, 229105823, 229105823,
              256670830, 256670830, 256670830, 256670830, 143639106, 143639106, 143639106, 143639106}))
  stage_6_butterfly_0 (
    .x_in(stage_5_per_out[0]),
    .y_in(stage_5_per_out[1]),
    .x_out(stage_6_per_in[0]),
    .y_out(stage_6_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 265190919, 265190919, 102773617, 102773617, 102773617, 102773617,
              210831626, 210831626, 210831626, 210831626, 84893967, 84893967, 84893967, 84893967,
              119480423, 119480423, 119480423, 119480423, 102579498, 102579498, 102579498, 102579498,
              129001811, 129001811, 129001811, 129001811, 72061017, 72061017, 72061017, 72061017,
              72052889, 72052889, 72052889, 72052889, 73825164, 73825164, 73825164, 73825164,
              18533839, 18533839, 18533839, 18533839, 168579404, 168579404, 168579404, 168579404,
              47877183, 47877183, 47877183, 47877183, 184798272, 184798272, 184798272, 184798272,
              5258704, 5258704, 5258704, 5258704, 92744225, 92744225, 92744225, 92744225,
              221840088, 221840088, 221840088, 221840088, 216372172, 216372172, 216372172, 216372172,
              231414272, 231414272, 231414272, 231414272, 94135184, 94135184, 94135184, 94135184,
              89995519, 89995519, 89995519, 89995519, 220656190, 220656190, 220656190, 220656190,
              183300662, 183300662, 183300662, 183300662, 160020761, 160020761, 160020761, 160020761,
              249274747, 249274747, 249274747, 249274747, 62061822, 62061822, 62061822, 62061822,
              76573097, 76573097, 76573097, 76573097, 35289455, 35289455, 35289455, 35289455,
              234642902, 234642902, 234642902, 234642902, 229105823, 229105823, 229105823, 229105823,
              256670830, 256670830, 256670830, 256670830, 143639106, 143639106, 143639106, 143639106}))
  stage_6_butterfly_1 (
    .x_in(stage_5_per_out[2]),
    .y_in(stage_5_per_out[3]),
    .x_out(stage_6_per_in[2]),
    .y_out(stage_6_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 265190919, 265190919, 102773617, 102773617, 102773617, 102773617,
              210831626, 210831626, 210831626, 210831626, 84893967, 84893967, 84893967, 84893967,
              119480423, 119480423, 119480423, 119480423, 102579498, 102579498, 102579498, 102579498,
              129001811, 129001811, 129001811, 129001811, 72061017, 72061017, 72061017, 72061017,
              72052889, 72052889, 72052889, 72052889, 73825164, 73825164, 73825164, 73825164,
              18533839, 18533839, 18533839, 18533839, 168579404, 168579404, 168579404, 168579404,
              47877183, 47877183, 47877183, 47877183, 184798272, 184798272, 184798272, 184798272,
              5258704, 5258704, 5258704, 5258704, 92744225, 92744225, 92744225, 92744225,
              221840088, 221840088, 221840088, 221840088, 216372172, 216372172, 216372172, 216372172,
              231414272, 231414272, 231414272, 231414272, 94135184, 94135184, 94135184, 94135184,
              89995519, 89995519, 89995519, 89995519, 220656190, 220656190, 220656190, 220656190,
              183300662, 183300662, 183300662, 183300662, 160020761, 160020761, 160020761, 160020761,
              249274747, 249274747, 249274747, 249274747, 62061822, 62061822, 62061822, 62061822,
              76573097, 76573097, 76573097, 76573097, 35289455, 35289455, 35289455, 35289455,
              234642902, 234642902, 234642902, 234642902, 229105823, 229105823, 229105823, 229105823,
              256670830, 256670830, 256670830, 256670830, 143639106, 143639106, 143639106, 143639106}))
  stage_6_butterfly_2 (
    .x_in(stage_5_per_out[4]),
    .y_in(stage_5_per_out[5]),
    .x_out(stage_6_per_in[4]),
    .y_out(stage_6_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 265190919, 265190919, 102773617, 102773617, 102773617, 102773617,
              210831626, 210831626, 210831626, 210831626, 84893967, 84893967, 84893967, 84893967,
              119480423, 119480423, 119480423, 119480423, 102579498, 102579498, 102579498, 102579498,
              129001811, 129001811, 129001811, 129001811, 72061017, 72061017, 72061017, 72061017,
              72052889, 72052889, 72052889, 72052889, 73825164, 73825164, 73825164, 73825164,
              18533839, 18533839, 18533839, 18533839, 168579404, 168579404, 168579404, 168579404,
              47877183, 47877183, 47877183, 47877183, 184798272, 184798272, 184798272, 184798272,
              5258704, 5258704, 5258704, 5258704, 92744225, 92744225, 92744225, 92744225,
              221840088, 221840088, 221840088, 221840088, 216372172, 216372172, 216372172, 216372172,
              231414272, 231414272, 231414272, 231414272, 94135184, 94135184, 94135184, 94135184,
              89995519, 89995519, 89995519, 89995519, 220656190, 220656190, 220656190, 220656190,
              183300662, 183300662, 183300662, 183300662, 160020761, 160020761, 160020761, 160020761,
              249274747, 249274747, 249274747, 249274747, 62061822, 62061822, 62061822, 62061822,
              76573097, 76573097, 76573097, 76573097, 35289455, 35289455, 35289455, 35289455,
              234642902, 234642902, 234642902, 234642902, 229105823, 229105823, 229105823, 229105823,
              256670830, 256670830, 256670830, 256670830, 143639106, 143639106, 143639106, 143639106}))
  stage_6_butterfly_3 (
    .x_in(stage_5_per_out[6]),
    .y_in(stage_5_per_out[7]),
    .x_out(stage_6_per_in[6]),
    .y_out(stage_6_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 265190919, 265190919, 102773617, 102773617, 102773617, 102773617,
              210831626, 210831626, 210831626, 210831626, 84893967, 84893967, 84893967, 84893967,
              119480423, 119480423, 119480423, 119480423, 102579498, 102579498, 102579498, 102579498,
              129001811, 129001811, 129001811, 129001811, 72061017, 72061017, 72061017, 72061017,
              72052889, 72052889, 72052889, 72052889, 73825164, 73825164, 73825164, 73825164,
              18533839, 18533839, 18533839, 18533839, 168579404, 168579404, 168579404, 168579404,
              47877183, 47877183, 47877183, 47877183, 184798272, 184798272, 184798272, 184798272,
              5258704, 5258704, 5258704, 5258704, 92744225, 92744225, 92744225, 92744225,
              221840088, 221840088, 221840088, 221840088, 216372172, 216372172, 216372172, 216372172,
              231414272, 231414272, 231414272, 231414272, 94135184, 94135184, 94135184, 94135184,
              89995519, 89995519, 89995519, 89995519, 220656190, 220656190, 220656190, 220656190,
              183300662, 183300662, 183300662, 183300662, 160020761, 160020761, 160020761, 160020761,
              249274747, 249274747, 249274747, 249274747, 62061822, 62061822, 62061822, 62061822,
              76573097, 76573097, 76573097, 76573097, 35289455, 35289455, 35289455, 35289455,
              234642902, 234642902, 234642902, 234642902, 229105823, 229105823, 229105823, 229105823,
              256670830, 256670830, 256670830, 256670830, 143639106, 143639106, 143639106, 143639106}))
  stage_6_butterfly_4 (
    .x_in(stage_5_per_out[8]),
    .y_in(stage_5_per_out[9]),
    .x_out(stage_6_per_in[8]),
    .y_out(stage_6_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 265190919, 265190919, 102773617, 102773617, 102773617, 102773617,
              210831626, 210831626, 210831626, 210831626, 84893967, 84893967, 84893967, 84893967,
              119480423, 119480423, 119480423, 119480423, 102579498, 102579498, 102579498, 102579498,
              129001811, 129001811, 129001811, 129001811, 72061017, 72061017, 72061017, 72061017,
              72052889, 72052889, 72052889, 72052889, 73825164, 73825164, 73825164, 73825164,
              18533839, 18533839, 18533839, 18533839, 168579404, 168579404, 168579404, 168579404,
              47877183, 47877183, 47877183, 47877183, 184798272, 184798272, 184798272, 184798272,
              5258704, 5258704, 5258704, 5258704, 92744225, 92744225, 92744225, 92744225,
              221840088, 221840088, 221840088, 221840088, 216372172, 216372172, 216372172, 216372172,
              231414272, 231414272, 231414272, 231414272, 94135184, 94135184, 94135184, 94135184,
              89995519, 89995519, 89995519, 89995519, 220656190, 220656190, 220656190, 220656190,
              183300662, 183300662, 183300662, 183300662, 160020761, 160020761, 160020761, 160020761,
              249274747, 249274747, 249274747, 249274747, 62061822, 62061822, 62061822, 62061822,
              76573097, 76573097, 76573097, 76573097, 35289455, 35289455, 35289455, 35289455,
              234642902, 234642902, 234642902, 234642902, 229105823, 229105823, 229105823, 229105823,
              256670830, 256670830, 256670830, 256670830, 143639106, 143639106, 143639106, 143639106}))
  stage_6_butterfly_5 (
    .x_in(stage_5_per_out[10]),
    .y_in(stage_5_per_out[11]),
    .x_out(stage_6_per_in[10]),
    .y_out(stage_6_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 265190919, 265190919, 102773617, 102773617, 102773617, 102773617,
              210831626, 210831626, 210831626, 210831626, 84893967, 84893967, 84893967, 84893967,
              119480423, 119480423, 119480423, 119480423, 102579498, 102579498, 102579498, 102579498,
              129001811, 129001811, 129001811, 129001811, 72061017, 72061017, 72061017, 72061017,
              72052889, 72052889, 72052889, 72052889, 73825164, 73825164, 73825164, 73825164,
              18533839, 18533839, 18533839, 18533839, 168579404, 168579404, 168579404, 168579404,
              47877183, 47877183, 47877183, 47877183, 184798272, 184798272, 184798272, 184798272,
              5258704, 5258704, 5258704, 5258704, 92744225, 92744225, 92744225, 92744225,
              221840088, 221840088, 221840088, 221840088, 216372172, 216372172, 216372172, 216372172,
              231414272, 231414272, 231414272, 231414272, 94135184, 94135184, 94135184, 94135184,
              89995519, 89995519, 89995519, 89995519, 220656190, 220656190, 220656190, 220656190,
              183300662, 183300662, 183300662, 183300662, 160020761, 160020761, 160020761, 160020761,
              249274747, 249274747, 249274747, 249274747, 62061822, 62061822, 62061822, 62061822,
              76573097, 76573097, 76573097, 76573097, 35289455, 35289455, 35289455, 35289455,
              234642902, 234642902, 234642902, 234642902, 229105823, 229105823, 229105823, 229105823,
              256670830, 256670830, 256670830, 256670830, 143639106, 143639106, 143639106, 143639106}))
  stage_6_butterfly_6 (
    .x_in(stage_5_per_out[12]),
    .y_in(stage_5_per_out[13]),
    .x_out(stage_6_per_in[12]),
    .y_out(stage_6_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 265190919, 265190919, 102773617, 102773617, 102773617, 102773617,
              210831626, 210831626, 210831626, 210831626, 84893967, 84893967, 84893967, 84893967,
              119480423, 119480423, 119480423, 119480423, 102579498, 102579498, 102579498, 102579498,
              129001811, 129001811, 129001811, 129001811, 72061017, 72061017, 72061017, 72061017,
              72052889, 72052889, 72052889, 72052889, 73825164, 73825164, 73825164, 73825164,
              18533839, 18533839, 18533839, 18533839, 168579404, 168579404, 168579404, 168579404,
              47877183, 47877183, 47877183, 47877183, 184798272, 184798272, 184798272, 184798272,
              5258704, 5258704, 5258704, 5258704, 92744225, 92744225, 92744225, 92744225,
              221840088, 221840088, 221840088, 221840088, 216372172, 216372172, 216372172, 216372172,
              231414272, 231414272, 231414272, 231414272, 94135184, 94135184, 94135184, 94135184,
              89995519, 89995519, 89995519, 89995519, 220656190, 220656190, 220656190, 220656190,
              183300662, 183300662, 183300662, 183300662, 160020761, 160020761, 160020761, 160020761,
              249274747, 249274747, 249274747, 249274747, 62061822, 62061822, 62061822, 62061822,
              76573097, 76573097, 76573097, 76573097, 35289455, 35289455, 35289455, 35289455,
              234642902, 234642902, 234642902, 234642902, 229105823, 229105823, 229105823, 229105823,
              256670830, 256670830, 256670830, 256670830, 143639106, 143639106, 143639106, 143639106}))
  stage_6_butterfly_7 (
    .x_in(stage_5_per_out[14]),
    .y_in(stage_5_per_out[15]),
    .x_out(stage_6_per_in[14]),
    .y_out(stage_6_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 265190919, 265190919, 102773617, 102773617, 102773617, 102773617,
              210831626, 210831626, 210831626, 210831626, 84893967, 84893967, 84893967, 84893967,
              119480423, 119480423, 119480423, 119480423, 102579498, 102579498, 102579498, 102579498,
              129001811, 129001811, 129001811, 129001811, 72061017, 72061017, 72061017, 72061017,
              72052889, 72052889, 72052889, 72052889, 73825164, 73825164, 73825164, 73825164,
              18533839, 18533839, 18533839, 18533839, 168579404, 168579404, 168579404, 168579404,
              47877183, 47877183, 47877183, 47877183, 184798272, 184798272, 184798272, 184798272,
              5258704, 5258704, 5258704, 5258704, 92744225, 92744225, 92744225, 92744225,
              221840088, 221840088, 221840088, 221840088, 216372172, 216372172, 216372172, 216372172,
              231414272, 231414272, 231414272, 231414272, 94135184, 94135184, 94135184, 94135184,
              89995519, 89995519, 89995519, 89995519, 220656190, 220656190, 220656190, 220656190,
              183300662, 183300662, 183300662, 183300662, 160020761, 160020761, 160020761, 160020761,
              249274747, 249274747, 249274747, 249274747, 62061822, 62061822, 62061822, 62061822,
              76573097, 76573097, 76573097, 76573097, 35289455, 35289455, 35289455, 35289455,
              234642902, 234642902, 234642902, 234642902, 229105823, 229105823, 229105823, 229105823,
              256670830, 256670830, 256670830, 256670830, 143639106, 143639106, 143639106, 143639106}))
  stage_6_butterfly_8 (
    .x_in(stage_5_per_out[16]),
    .y_in(stage_5_per_out[17]),
    .x_out(stage_6_per_in[16]),
    .y_out(stage_6_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 265190919, 265190919, 102773617, 102773617, 102773617, 102773617,
              210831626, 210831626, 210831626, 210831626, 84893967, 84893967, 84893967, 84893967,
              119480423, 119480423, 119480423, 119480423, 102579498, 102579498, 102579498, 102579498,
              129001811, 129001811, 129001811, 129001811, 72061017, 72061017, 72061017, 72061017,
              72052889, 72052889, 72052889, 72052889, 73825164, 73825164, 73825164, 73825164,
              18533839, 18533839, 18533839, 18533839, 168579404, 168579404, 168579404, 168579404,
              47877183, 47877183, 47877183, 47877183, 184798272, 184798272, 184798272, 184798272,
              5258704, 5258704, 5258704, 5258704, 92744225, 92744225, 92744225, 92744225,
              221840088, 221840088, 221840088, 221840088, 216372172, 216372172, 216372172, 216372172,
              231414272, 231414272, 231414272, 231414272, 94135184, 94135184, 94135184, 94135184,
              89995519, 89995519, 89995519, 89995519, 220656190, 220656190, 220656190, 220656190,
              183300662, 183300662, 183300662, 183300662, 160020761, 160020761, 160020761, 160020761,
              249274747, 249274747, 249274747, 249274747, 62061822, 62061822, 62061822, 62061822,
              76573097, 76573097, 76573097, 76573097, 35289455, 35289455, 35289455, 35289455,
              234642902, 234642902, 234642902, 234642902, 229105823, 229105823, 229105823, 229105823,
              256670830, 256670830, 256670830, 256670830, 143639106, 143639106, 143639106, 143639106}))
  stage_6_butterfly_9 (
    .x_in(stage_5_per_out[18]),
    .y_in(stage_5_per_out[19]),
    .x_out(stage_6_per_in[18]),
    .y_out(stage_6_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 265190919, 265190919, 102773617, 102773617, 102773617, 102773617,
              210831626, 210831626, 210831626, 210831626, 84893967, 84893967, 84893967, 84893967,
              119480423, 119480423, 119480423, 119480423, 102579498, 102579498, 102579498, 102579498,
              129001811, 129001811, 129001811, 129001811, 72061017, 72061017, 72061017, 72061017,
              72052889, 72052889, 72052889, 72052889, 73825164, 73825164, 73825164, 73825164,
              18533839, 18533839, 18533839, 18533839, 168579404, 168579404, 168579404, 168579404,
              47877183, 47877183, 47877183, 47877183, 184798272, 184798272, 184798272, 184798272,
              5258704, 5258704, 5258704, 5258704, 92744225, 92744225, 92744225, 92744225,
              221840088, 221840088, 221840088, 221840088, 216372172, 216372172, 216372172, 216372172,
              231414272, 231414272, 231414272, 231414272, 94135184, 94135184, 94135184, 94135184,
              89995519, 89995519, 89995519, 89995519, 220656190, 220656190, 220656190, 220656190,
              183300662, 183300662, 183300662, 183300662, 160020761, 160020761, 160020761, 160020761,
              249274747, 249274747, 249274747, 249274747, 62061822, 62061822, 62061822, 62061822,
              76573097, 76573097, 76573097, 76573097, 35289455, 35289455, 35289455, 35289455,
              234642902, 234642902, 234642902, 234642902, 229105823, 229105823, 229105823, 229105823,
              256670830, 256670830, 256670830, 256670830, 143639106, 143639106, 143639106, 143639106}))
  stage_6_butterfly_10 (
    .x_in(stage_5_per_out[20]),
    .y_in(stage_5_per_out[21]),
    .x_out(stage_6_per_in[20]),
    .y_out(stage_6_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 265190919, 265190919, 102773617, 102773617, 102773617, 102773617,
              210831626, 210831626, 210831626, 210831626, 84893967, 84893967, 84893967, 84893967,
              119480423, 119480423, 119480423, 119480423, 102579498, 102579498, 102579498, 102579498,
              129001811, 129001811, 129001811, 129001811, 72061017, 72061017, 72061017, 72061017,
              72052889, 72052889, 72052889, 72052889, 73825164, 73825164, 73825164, 73825164,
              18533839, 18533839, 18533839, 18533839, 168579404, 168579404, 168579404, 168579404,
              47877183, 47877183, 47877183, 47877183, 184798272, 184798272, 184798272, 184798272,
              5258704, 5258704, 5258704, 5258704, 92744225, 92744225, 92744225, 92744225,
              221840088, 221840088, 221840088, 221840088, 216372172, 216372172, 216372172, 216372172,
              231414272, 231414272, 231414272, 231414272, 94135184, 94135184, 94135184, 94135184,
              89995519, 89995519, 89995519, 89995519, 220656190, 220656190, 220656190, 220656190,
              183300662, 183300662, 183300662, 183300662, 160020761, 160020761, 160020761, 160020761,
              249274747, 249274747, 249274747, 249274747, 62061822, 62061822, 62061822, 62061822,
              76573097, 76573097, 76573097, 76573097, 35289455, 35289455, 35289455, 35289455,
              234642902, 234642902, 234642902, 234642902, 229105823, 229105823, 229105823, 229105823,
              256670830, 256670830, 256670830, 256670830, 143639106, 143639106, 143639106, 143639106}))
  stage_6_butterfly_11 (
    .x_in(stage_5_per_out[22]),
    .y_in(stage_5_per_out[23]),
    .x_out(stage_6_per_in[22]),
    .y_out(stage_6_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 265190919, 265190919, 102773617, 102773617, 102773617, 102773617,
              210831626, 210831626, 210831626, 210831626, 84893967, 84893967, 84893967, 84893967,
              119480423, 119480423, 119480423, 119480423, 102579498, 102579498, 102579498, 102579498,
              129001811, 129001811, 129001811, 129001811, 72061017, 72061017, 72061017, 72061017,
              72052889, 72052889, 72052889, 72052889, 73825164, 73825164, 73825164, 73825164,
              18533839, 18533839, 18533839, 18533839, 168579404, 168579404, 168579404, 168579404,
              47877183, 47877183, 47877183, 47877183, 184798272, 184798272, 184798272, 184798272,
              5258704, 5258704, 5258704, 5258704, 92744225, 92744225, 92744225, 92744225,
              221840088, 221840088, 221840088, 221840088, 216372172, 216372172, 216372172, 216372172,
              231414272, 231414272, 231414272, 231414272, 94135184, 94135184, 94135184, 94135184,
              89995519, 89995519, 89995519, 89995519, 220656190, 220656190, 220656190, 220656190,
              183300662, 183300662, 183300662, 183300662, 160020761, 160020761, 160020761, 160020761,
              249274747, 249274747, 249274747, 249274747, 62061822, 62061822, 62061822, 62061822,
              76573097, 76573097, 76573097, 76573097, 35289455, 35289455, 35289455, 35289455,
              234642902, 234642902, 234642902, 234642902, 229105823, 229105823, 229105823, 229105823,
              256670830, 256670830, 256670830, 256670830, 143639106, 143639106, 143639106, 143639106}))
  stage_6_butterfly_12 (
    .x_in(stage_5_per_out[24]),
    .y_in(stage_5_per_out[25]),
    .x_out(stage_6_per_in[24]),
    .y_out(stage_6_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 265190919, 265190919, 102773617, 102773617, 102773617, 102773617,
              210831626, 210831626, 210831626, 210831626, 84893967, 84893967, 84893967, 84893967,
              119480423, 119480423, 119480423, 119480423, 102579498, 102579498, 102579498, 102579498,
              129001811, 129001811, 129001811, 129001811, 72061017, 72061017, 72061017, 72061017,
              72052889, 72052889, 72052889, 72052889, 73825164, 73825164, 73825164, 73825164,
              18533839, 18533839, 18533839, 18533839, 168579404, 168579404, 168579404, 168579404,
              47877183, 47877183, 47877183, 47877183, 184798272, 184798272, 184798272, 184798272,
              5258704, 5258704, 5258704, 5258704, 92744225, 92744225, 92744225, 92744225,
              221840088, 221840088, 221840088, 221840088, 216372172, 216372172, 216372172, 216372172,
              231414272, 231414272, 231414272, 231414272, 94135184, 94135184, 94135184, 94135184,
              89995519, 89995519, 89995519, 89995519, 220656190, 220656190, 220656190, 220656190,
              183300662, 183300662, 183300662, 183300662, 160020761, 160020761, 160020761, 160020761,
              249274747, 249274747, 249274747, 249274747, 62061822, 62061822, 62061822, 62061822,
              76573097, 76573097, 76573097, 76573097, 35289455, 35289455, 35289455, 35289455,
              234642902, 234642902, 234642902, 234642902, 229105823, 229105823, 229105823, 229105823,
              256670830, 256670830, 256670830, 256670830, 143639106, 143639106, 143639106, 143639106}))
  stage_6_butterfly_13 (
    .x_in(stage_5_per_out[26]),
    .y_in(stage_5_per_out[27]),
    .x_out(stage_6_per_in[26]),
    .y_out(stage_6_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 265190919, 265190919, 102773617, 102773617, 102773617, 102773617,
              210831626, 210831626, 210831626, 210831626, 84893967, 84893967, 84893967, 84893967,
              119480423, 119480423, 119480423, 119480423, 102579498, 102579498, 102579498, 102579498,
              129001811, 129001811, 129001811, 129001811, 72061017, 72061017, 72061017, 72061017,
              72052889, 72052889, 72052889, 72052889, 73825164, 73825164, 73825164, 73825164,
              18533839, 18533839, 18533839, 18533839, 168579404, 168579404, 168579404, 168579404,
              47877183, 47877183, 47877183, 47877183, 184798272, 184798272, 184798272, 184798272,
              5258704, 5258704, 5258704, 5258704, 92744225, 92744225, 92744225, 92744225,
              221840088, 221840088, 221840088, 221840088, 216372172, 216372172, 216372172, 216372172,
              231414272, 231414272, 231414272, 231414272, 94135184, 94135184, 94135184, 94135184,
              89995519, 89995519, 89995519, 89995519, 220656190, 220656190, 220656190, 220656190,
              183300662, 183300662, 183300662, 183300662, 160020761, 160020761, 160020761, 160020761,
              249274747, 249274747, 249274747, 249274747, 62061822, 62061822, 62061822, 62061822,
              76573097, 76573097, 76573097, 76573097, 35289455, 35289455, 35289455, 35289455,
              234642902, 234642902, 234642902, 234642902, 229105823, 229105823, 229105823, 229105823,
              256670830, 256670830, 256670830, 256670830, 143639106, 143639106, 143639106, 143639106}))
  stage_6_butterfly_14 (
    .x_in(stage_5_per_out[28]),
    .y_in(stage_5_per_out[29]),
    .x_out(stage_6_per_in[28]),
    .y_out(stage_6_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[6]),
    .factors({265190919, 265190919, 265190919, 265190919, 102773617, 102773617, 102773617, 102773617,
              210831626, 210831626, 210831626, 210831626, 84893967, 84893967, 84893967, 84893967,
              119480423, 119480423, 119480423, 119480423, 102579498, 102579498, 102579498, 102579498,
              129001811, 129001811, 129001811, 129001811, 72061017, 72061017, 72061017, 72061017,
              72052889, 72052889, 72052889, 72052889, 73825164, 73825164, 73825164, 73825164,
              18533839, 18533839, 18533839, 18533839, 168579404, 168579404, 168579404, 168579404,
              47877183, 47877183, 47877183, 47877183, 184798272, 184798272, 184798272, 184798272,
              5258704, 5258704, 5258704, 5258704, 92744225, 92744225, 92744225, 92744225,
              221840088, 221840088, 221840088, 221840088, 216372172, 216372172, 216372172, 216372172,
              231414272, 231414272, 231414272, 231414272, 94135184, 94135184, 94135184, 94135184,
              89995519, 89995519, 89995519, 89995519, 220656190, 220656190, 220656190, 220656190,
              183300662, 183300662, 183300662, 183300662, 160020761, 160020761, 160020761, 160020761,
              249274747, 249274747, 249274747, 249274747, 62061822, 62061822, 62061822, 62061822,
              76573097, 76573097, 76573097, 76573097, 35289455, 35289455, 35289455, 35289455,
              234642902, 234642902, 234642902, 234642902, 229105823, 229105823, 229105823, 229105823,
              256670830, 256670830, 256670830, 256670830, 143639106, 143639106, 143639106, 143639106}))
  stage_6_butterfly_15 (
    .x_in(stage_5_per_out[30]),
    .y_in(stage_5_per_out[31]),
    .x_out(stage_6_per_in[30]),
    .y_out(stage_6_per_in[31]),
    .clk(clk),
    .rst(rst)
  );






  // TODO(Yang): stage 6 -> stage 7 permutation
  // FIXME: ignore butterfly units for now.
  stage_6_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_6_7_per (
    .inData_0(stage_6_per_in[0]),
    .inData_1(stage_6_per_in[1]),
    .inData_2(stage_6_per_in[2]),
    .inData_3(stage_6_per_in[3]),
    .inData_4(stage_6_per_in[4]),
    .inData_5(stage_6_per_in[5]),
    .inData_6(stage_6_per_in[6]),
    .inData_7(stage_6_per_in[7]),
    .inData_8(stage_6_per_in[8]),
    .inData_9(stage_6_per_in[9]),
    .inData_10(stage_6_per_in[10]),
    .inData_11(stage_6_per_in[11]),
    .inData_12(stage_6_per_in[12]),
    .inData_13(stage_6_per_in[13]),
    .inData_14(stage_6_per_in[14]),
    .inData_15(stage_6_per_in[15]),
    .inData_16(stage_6_per_in[16]),
    .inData_17(stage_6_per_in[17]),
    .inData_18(stage_6_per_in[18]),
    .inData_19(stage_6_per_in[19]),
    .inData_20(stage_6_per_in[20]),
    .inData_21(stage_6_per_in[21]),
    .inData_22(stage_6_per_in[22]),
    .inData_23(stage_6_per_in[23]),
    .inData_24(stage_6_per_in[24]),
    .inData_25(stage_6_per_in[25]),
    .inData_26(stage_6_per_in[26]),
    .inData_27(stage_6_per_in[27]),
    .inData_28(stage_6_per_in[28]),
    .inData_29(stage_6_per_in[29]),
    .inData_30(stage_6_per_in[30]),
    .inData_31(stage_6_per_in[31]),
    .outData_0(stage_6_per_out[0]),
    .outData_1(stage_6_per_out[1]),
    .outData_2(stage_6_per_out[2]),
    .outData_3(stage_6_per_out[3]),
    .outData_4(stage_6_per_out[4]),
    .outData_5(stage_6_per_out[5]),
    .outData_6(stage_6_per_out[6]),
    .outData_7(stage_6_per_out[7]),
    .outData_8(stage_6_per_out[8]),
    .outData_9(stage_6_per_out[9]),
    .outData_10(stage_6_per_out[10]),
    .outData_11(stage_6_per_out[11]),
    .outData_12(stage_6_per_out[12]),
    .outData_13(stage_6_per_out[13]),
    .outData_14(stage_6_per_out[14]),
    .outData_15(stage_6_per_out[15]),
    .outData_16(stage_6_per_out[16]),
    .outData_17(stage_6_per_out[17]),
    .outData_18(stage_6_per_out[18]),
    .outData_19(stage_6_per_out[19]),
    .outData_20(stage_6_per_out[20]),
    .outData_21(stage_6_per_out[21]),
    .outData_22(stage_6_per_out[22]),
    .outData_23(stage_6_per_out[23]),
    .outData_24(stage_6_per_out[24]),
    .outData_25(stage_6_per_out[25]),
    .outData_26(stage_6_per_out[26]),
    .outData_27(stage_6_per_out[27]),
    .outData_28(stage_6_per_out[28]),
    .outData_29(stage_6_per_out[29]),
    .outData_30(stage_6_per_out[30]),
    .outData_31(stage_6_per_out[31]),
    .in_start(in_start[6]),
    .out_start(out_start[6]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 7 32 butterfly units
  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907,
              33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015,
              69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111,
              155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162,
              57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932,
              225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267,
              73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048,
              25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445,
              70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_0 (
    .x_in(stage_6_per_out[0]),
    .y_in(stage_6_per_out[1]),
    .x_out(stage_7_per_in[0]),
    .y_out(stage_7_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907,
              33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015,
              69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111,
              155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162,
              57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932,
              225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267,
              73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048,
              25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445,
              70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_1 (
    .x_in(stage_6_per_out[2]),
    .y_in(stage_6_per_out[3]),
    .x_out(stage_7_per_in[2]),
    .y_out(stage_7_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907,
              33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015,
              69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111,
              155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162,
              57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932,
              225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267,
              73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048,
              25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445,
              70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_2 (
    .x_in(stage_6_per_out[4]),
    .y_in(stage_6_per_out[5]),
    .x_out(stage_7_per_in[4]),
    .y_out(stage_7_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907,
              33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015,
              69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111,
              155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162,
              57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932,
              225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267,
              73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048,
              25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445,
              70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_3 (
    .x_in(stage_6_per_out[6]),
    .y_in(stage_6_per_out[7]),
    .x_out(stage_7_per_in[6]),
    .y_out(stage_7_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907,
              33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015,
              69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111,
              155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162,
              57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932,
              225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267,
              73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048,
              25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445,
              70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_4 (
    .x_in(stage_6_per_out[8]),
    .y_in(stage_6_per_out[9]),
    .x_out(stage_7_per_in[8]),
    .y_out(stage_7_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907,
              33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015,
              69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111,
              155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162,
              57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932,
              225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267,
              73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048,
              25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445,
              70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_5 (
    .x_in(stage_6_per_out[10]),
    .y_in(stage_6_per_out[11]),
    .x_out(stage_7_per_in[10]),
    .y_out(stage_7_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907,
              33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015,
              69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111,
              155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162,
              57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932,
              225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267,
              73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048,
              25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445,
              70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_6 (
    .x_in(stage_6_per_out[12]),
    .y_in(stage_6_per_out[13]),
    .x_out(stage_7_per_in[12]),
    .y_out(stage_7_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907,
              33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015,
              69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111,
              155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162,
              57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932,
              225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267,
              73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048,
              25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445,
              70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_7 (
    .x_in(stage_6_per_out[14]),
    .y_in(stage_6_per_out[15]),
    .x_out(stage_7_per_in[14]),
    .y_out(stage_7_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907,
              33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015,
              69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111,
              155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162,
              57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932,
              225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267,
              73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048,
              25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445,
              70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_8 (
    .x_in(stage_6_per_out[16]),
    .y_in(stage_6_per_out[17]),
    .x_out(stage_7_per_in[16]),
    .y_out(stage_7_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907,
              33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015,
              69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111,
              155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162,
              57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932,
              225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267,
              73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048,
              25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445,
              70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_9 (
    .x_in(stage_6_per_out[18]),
    .y_in(stage_6_per_out[19]),
    .x_out(stage_7_per_in[18]),
    .y_out(stage_7_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907,
              33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015,
              69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111,
              155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162,
              57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932,
              225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267,
              73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048,
              25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445,
              70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_10 (
    .x_in(stage_6_per_out[20]),
    .y_in(stage_6_per_out[21]),
    .x_out(stage_7_per_in[20]),
    .y_out(stage_7_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907,
              33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015,
              69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111,
              155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162,
              57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932,
              225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267,
              73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048,
              25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445,
              70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_11 (
    .x_in(stage_6_per_out[22]),
    .y_in(stage_6_per_out[23]),
    .x_out(stage_7_per_in[22]),
    .y_out(stage_7_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907,
              33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015,
              69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111,
              155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162,
              57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932,
              225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267,
              73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048,
              25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445,
              70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_12 (
    .x_in(stage_6_per_out[24]),
    .y_in(stage_6_per_out[25]),
    .x_out(stage_7_per_in[24]),
    .y_out(stage_7_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907,
              33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015,
              69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111,
              155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162,
              57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932,
              225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267,
              73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048,
              25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445,
              70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_13 (
    .x_in(stage_6_per_out[26]),
    .y_in(stage_6_per_out[27]),
    .x_out(stage_7_per_in[26]),
    .y_out(stage_7_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907,
              33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015,
              69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111,
              155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162,
              57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932,
              225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267,
              73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048,
              25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445,
              70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_14 (
    .x_in(stage_6_per_out[28]),
    .y_in(stage_6_per_out[29]),
    .x_out(stage_7_per_in[28]),
    .y_out(stage_7_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[7]),
    .factors({47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907, 47600907,
              33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981, 33383981,
              125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015, 125976015,
              69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086, 69075086,
              7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111, 7802111,
              155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840, 155624840,
              134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162, 134587162,
              57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092, 57620092,
              133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932, 133035932,
              225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856, 225387856,
              163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267, 163057267,
              73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196, 73648196,
              46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048, 46265048,
              25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822, 25800822,
              136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445, 136955445,
              70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281, 70516281}))
  stage_7_butterfly_15 (
    .x_in(stage_6_per_out[30]),
    .y_in(stage_6_per_out[31]),
    .x_out(stage_7_per_in[30]),
    .y_out(stage_7_per_in[31]),
    .clk(clk),
    .rst(rst)
  );






  // TODO(Yang): stage 7 -> stage 8 permutation
  // FIXME: ignore butterfly units for now.
  stage_7_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_7_8_per (
    .inData_0(stage_7_per_in[0]),
    .inData_1(stage_7_per_in[1]),
    .inData_2(stage_7_per_in[2]),
    .inData_3(stage_7_per_in[3]),
    .inData_4(stage_7_per_in[4]),
    .inData_5(stage_7_per_in[5]),
    .inData_6(stage_7_per_in[6]),
    .inData_7(stage_7_per_in[7]),
    .inData_8(stage_7_per_in[8]),
    .inData_9(stage_7_per_in[9]),
    .inData_10(stage_7_per_in[10]),
    .inData_11(stage_7_per_in[11]),
    .inData_12(stage_7_per_in[12]),
    .inData_13(stage_7_per_in[13]),
    .inData_14(stage_7_per_in[14]),
    .inData_15(stage_7_per_in[15]),
    .inData_16(stage_7_per_in[16]),
    .inData_17(stage_7_per_in[17]),
    .inData_18(stage_7_per_in[18]),
    .inData_19(stage_7_per_in[19]),
    .inData_20(stage_7_per_in[20]),
    .inData_21(stage_7_per_in[21]),
    .inData_22(stage_7_per_in[22]),
    .inData_23(stage_7_per_in[23]),
    .inData_24(stage_7_per_in[24]),
    .inData_25(stage_7_per_in[25]),
    .inData_26(stage_7_per_in[26]),
    .inData_27(stage_7_per_in[27]),
    .inData_28(stage_7_per_in[28]),
    .inData_29(stage_7_per_in[29]),
    .inData_30(stage_7_per_in[30]),
    .inData_31(stage_7_per_in[31]),
    .outData_0(stage_7_per_out[0]),
    .outData_1(stage_7_per_out[1]),
    .outData_2(stage_7_per_out[2]),
    .outData_3(stage_7_per_out[3]),
    .outData_4(stage_7_per_out[4]),
    .outData_5(stage_7_per_out[5]),
    .outData_6(stage_7_per_out[6]),
    .outData_7(stage_7_per_out[7]),
    .outData_8(stage_7_per_out[8]),
    .outData_9(stage_7_per_out[9]),
    .outData_10(stage_7_per_out[10]),
    .outData_11(stage_7_per_out[11]),
    .outData_12(stage_7_per_out[12]),
    .outData_13(stage_7_per_out[13]),
    .outData_14(stage_7_per_out[14]),
    .outData_15(stage_7_per_out[15]),
    .outData_16(stage_7_per_out[16]),
    .outData_17(stage_7_per_out[17]),
    .outData_18(stage_7_per_out[18]),
    .outData_19(stage_7_per_out[19]),
    .outData_20(stage_7_per_out[20]),
    .outData_21(stage_7_per_out[21]),
    .outData_22(stage_7_per_out[22]),
    .outData_23(stage_7_per_out[23]),
    .outData_24(stage_7_per_out[24]),
    .outData_25(stage_7_per_out[25]),
    .outData_26(stage_7_per_out[26]),
    .outData_27(stage_7_per_out[27]),
    .outData_28(stage_7_per_out[28]),
    .outData_29(stage_7_per_out[29]),
    .outData_30(stage_7_per_out[30]),
    .outData_31(stage_7_per_out[31]),
    .in_start(in_start[7]),
    .out_start(out_start[7]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 8 32 butterfly units
  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_0 (
    .x_in(stage_7_per_out[0]),
    .y_in(stage_7_per_out[1]),
    .x_out(stage_8_per_in[0]),
    .y_out(stage_8_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_1 (
    .x_in(stage_7_per_out[2]),
    .y_in(stage_7_per_out[3]),
    .x_out(stage_8_per_in[2]),
    .y_out(stage_8_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_2 (
    .x_in(stage_7_per_out[4]),
    .y_in(stage_7_per_out[5]),
    .x_out(stage_8_per_in[4]),
    .y_out(stage_8_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_3 (
    .x_in(stage_7_per_out[6]),
    .y_in(stage_7_per_out[7]),
    .x_out(stage_8_per_in[6]),
    .y_out(stage_8_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_4 (
    .x_in(stage_7_per_out[8]),
    .y_in(stage_7_per_out[9]),
    .x_out(stage_8_per_in[8]),
    .y_out(stage_8_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_5 (
    .x_in(stage_7_per_out[10]),
    .y_in(stage_7_per_out[11]),
    .x_out(stage_8_per_in[10]),
    .y_out(stage_8_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_6 (
    .x_in(stage_7_per_out[12]),
    .y_in(stage_7_per_out[13]),
    .x_out(stage_8_per_in[12]),
    .y_out(stage_8_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_7 (
    .x_in(stage_7_per_out[14]),
    .y_in(stage_7_per_out[15]),
    .x_out(stage_8_per_in[14]),
    .y_out(stage_8_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_8 (
    .x_in(stage_7_per_out[16]),
    .y_in(stage_7_per_out[17]),
    .x_out(stage_8_per_in[16]),
    .y_out(stage_8_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_9 (
    .x_in(stage_7_per_out[18]),
    .y_in(stage_7_per_out[19]),
    .x_out(stage_8_per_in[18]),
    .y_out(stage_8_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_10 (
    .x_in(stage_7_per_out[20]),
    .y_in(stage_7_per_out[21]),
    .x_out(stage_8_per_in[20]),
    .y_out(stage_8_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_11 (
    .x_in(stage_7_per_out[22]),
    .y_in(stage_7_per_out[23]),
    .x_out(stage_8_per_in[22]),
    .y_out(stage_8_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_12 (
    .x_in(stage_7_per_out[24]),
    .y_in(stage_7_per_out[25]),
    .x_out(stage_8_per_in[24]),
    .y_out(stage_8_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_13 (
    .x_in(stage_7_per_out[26]),
    .y_in(stage_7_per_out[27]),
    .x_out(stage_8_per_in[26]),
    .y_out(stage_8_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_14 (
    .x_in(stage_7_per_out[28]),
    .y_in(stage_7_per_out[29]),
    .x_out(stage_8_per_in[28]),
    .y_out(stage_8_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[8]),
    .factors({177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333, 177699333,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074, 105446074,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417, 197095417,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680, 140261680,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933, 87759933,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025, 172037025,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502, 48587502,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660,
              137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660, 137531660}))
  stage_8_butterfly_15 (
    .x_in(stage_7_per_out[30]),
    .y_in(stage_7_per_out[31]),
    .x_out(stage_8_per_in[30]),
    .y_out(stage_8_per_in[31]),
    .clk(clk),
    .rst(rst)
  );




  // TODO(Yang): stage 8 -> stage 9 permutation
  // FIXME: ignore butterfly units for now.
  stage_8_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_8_9_per (
    .inData_0(stage_8_per_in[0]),
    .inData_1(stage_8_per_in[1]),
    .inData_2(stage_8_per_in[2]),
    .inData_3(stage_8_per_in[3]),
    .inData_4(stage_8_per_in[4]),
    .inData_5(stage_8_per_in[5]),
    .inData_6(stage_8_per_in[6]),
    .inData_7(stage_8_per_in[7]),
    .inData_8(stage_8_per_in[8]),
    .inData_9(stage_8_per_in[9]),
    .inData_10(stage_8_per_in[10]),
    .inData_11(stage_8_per_in[11]),
    .inData_12(stage_8_per_in[12]),
    .inData_13(stage_8_per_in[13]),
    .inData_14(stage_8_per_in[14]),
    .inData_15(stage_8_per_in[15]),
    .inData_16(stage_8_per_in[16]),
    .inData_17(stage_8_per_in[17]),
    .inData_18(stage_8_per_in[18]),
    .inData_19(stage_8_per_in[19]),
    .inData_20(stage_8_per_in[20]),
    .inData_21(stage_8_per_in[21]),
    .inData_22(stage_8_per_in[22]),
    .inData_23(stage_8_per_in[23]),
    .inData_24(stage_8_per_in[24]),
    .inData_25(stage_8_per_in[25]),
    .inData_26(stage_8_per_in[26]),
    .inData_27(stage_8_per_in[27]),
    .inData_28(stage_8_per_in[28]),
    .inData_29(stage_8_per_in[29]),
    .inData_30(stage_8_per_in[30]),
    .inData_31(stage_8_per_in[31]),
    .outData_0(stage_8_per_out[0]),
    .outData_1(stage_8_per_out[1]),
    .outData_2(stage_8_per_out[2]),
    .outData_3(stage_8_per_out[3]),
    .outData_4(stage_8_per_out[4]),
    .outData_5(stage_8_per_out[5]),
    .outData_6(stage_8_per_out[6]),
    .outData_7(stage_8_per_out[7]),
    .outData_8(stage_8_per_out[8]),
    .outData_9(stage_8_per_out[9]),
    .outData_10(stage_8_per_out[10]),
    .outData_11(stage_8_per_out[11]),
    .outData_12(stage_8_per_out[12]),
    .outData_13(stage_8_per_out[13]),
    .outData_14(stage_8_per_out[14]),
    .outData_15(stage_8_per_out[15]),
    .outData_16(stage_8_per_out[16]),
    .outData_17(stage_8_per_out[17]),
    .outData_18(stage_8_per_out[18]),
    .outData_19(stage_8_per_out[19]),
    .outData_20(stage_8_per_out[20]),
    .outData_21(stage_8_per_out[21]),
    .outData_22(stage_8_per_out[22]),
    .outData_23(stage_8_per_out[23]),
    .outData_24(stage_8_per_out[24]),
    .outData_25(stage_8_per_out[25]),
    .outData_26(stage_8_per_out[26]),
    .outData_27(stage_8_per_out[27]),
    .outData_28(stage_8_per_out[28]),
    .outData_29(stage_8_per_out[29]),
    .outData_30(stage_8_per_out[30]),
    .outData_31(stage_8_per_out[31]),
    .in_start(in_start[8]),
    .out_start(out_start[8]),
    .clk(clk),
    .rst(rst)
  );
  // TODO(Tian): stage 9 32 butterfly units
  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_0 (
    .x_in(stage_8_per_out[0]),
    .y_in(stage_8_per_out[1]),
    .x_out(stage_9_per_in[0]),
    .y_out(stage_9_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_1 (
    .x_in(stage_8_per_out[2]),
    .y_in(stage_8_per_out[3]),
    .x_out(stage_9_per_in[2]),
    .y_out(stage_9_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_2 (
    .x_in(stage_8_per_out[4]),
    .y_in(stage_8_per_out[5]),
    .x_out(stage_9_per_in[4]),
    .y_out(stage_9_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_3 (
    .x_in(stage_8_per_out[6]),
    .y_in(stage_8_per_out[7]),
    .x_out(stage_9_per_in[6]),
    .y_out(stage_9_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_4 (
    .x_in(stage_8_per_out[8]),
    .y_in(stage_8_per_out[9]),
    .x_out(stage_9_per_in[8]),
    .y_out(stage_9_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_5 (
    .x_in(stage_8_per_out[10]),
    .y_in(stage_8_per_out[11]),
    .x_out(stage_9_per_in[10]),
    .y_out(stage_9_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_6 (
    .x_in(stage_8_per_out[12]),
    .y_in(stage_8_per_out[13]),
    .x_out(stage_9_per_in[12]),
    .y_out(stage_9_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_7 (
    .x_in(stage_8_per_out[14]),
    .y_in(stage_8_per_out[15]),
    .x_out(stage_9_per_in[14]),
    .y_out(stage_9_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_8 (
    .x_in(stage_8_per_out[16]),
    .y_in(stage_8_per_out[17]),
    .x_out(stage_9_per_in[16]),
    .y_out(stage_9_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_9 (
    .x_in(stage_8_per_out[18]),
    .y_in(stage_8_per_out[19]),
    .x_out(stage_9_per_in[18]),
    .y_out(stage_9_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_10 (
    .x_in(stage_8_per_out[20]),
    .y_in(stage_8_per_out[21]),
    .x_out(stage_9_per_in[20]),
    .y_out(stage_9_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_11 (
    .x_in(stage_8_per_out[22]),
    .y_in(stage_8_per_out[23]),
    .x_out(stage_9_per_in[22]),
    .y_out(stage_9_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_12 (
    .x_in(stage_8_per_out[24]),
    .y_in(stage_8_per_out[25]),
    .x_out(stage_9_per_in[24]),
    .y_out(stage_9_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_13 (
    .x_in(stage_8_per_out[26]),
    .y_in(stage_8_per_out[27]),
    .x_out(stage_9_per_in[26]),
    .y_out(stage_9_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_14 (
    .x_in(stage_8_per_out[28]),
    .y_in(stage_8_per_out[29]),
    .x_out(stage_9_per_in[28]),
    .y_out(stage_9_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[9]),
    .factors({198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595, 198795595,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716, 174860716,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461, 250183461,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115,
              88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115, 88202115}))
  stage_9_butterfly_15 (
    .x_in(stage_8_per_out[30]),
    .y_in(stage_8_per_out[31]),
    .x_out(stage_9_per_in[30]),
    .y_out(stage_9_per_in[31]),
    .clk(clk),
    .rst(rst)
  );


  // TODO(Yang): Update stride
  stage_9_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_9_10_per (
    .inData_0(stage_9_per_in[0]),
    .inData_1(stage_9_per_in[1]),
    .inData_2(stage_9_per_in[2]),
    .inData_3(stage_9_per_in[3]),
    .inData_4(stage_9_per_in[4]),
    .inData_5(stage_9_per_in[5]),
    .inData_6(stage_9_per_in[6]),
    .inData_7(stage_9_per_in[7]),
    .inData_8(stage_9_per_in[8]),
    .inData_9(stage_9_per_in[9]),
    .inData_10(stage_9_per_in[10]),
    .inData_11(stage_9_per_in[11]),
    .inData_12(stage_9_per_in[12]),
    .inData_13(stage_9_per_in[13]),
    .inData_14(stage_9_per_in[14]),
    .inData_15(stage_9_per_in[15]),
    .inData_16(stage_9_per_in[16]),
    .inData_17(stage_9_per_in[17]),
    .inData_18(stage_9_per_in[18]),
    .inData_19(stage_9_per_in[19]),
    .inData_20(stage_9_per_in[20]),
    .inData_21(stage_9_per_in[21]),
    .inData_22(stage_9_per_in[22]),
    .inData_23(stage_9_per_in[23]),
    .inData_24(stage_9_per_in[24]),
    .inData_25(stage_9_per_in[25]),
    .inData_26(stage_9_per_in[26]),
    .inData_27(stage_9_per_in[27]),
    .inData_28(stage_9_per_in[28]),
    .inData_29(stage_9_per_in[29]),
    .inData_30(stage_9_per_in[30]),
    .inData_31(stage_9_per_in[31]),
    .outData_0(stage_9_per_out[0]),
    .outData_1(stage_9_per_out[1]),
    .outData_2(stage_9_per_out[2]),
    .outData_3(stage_9_per_out[3]),
    .outData_4(stage_9_per_out[4]),
    .outData_5(stage_9_per_out[5]),
    .outData_6(stage_9_per_out[6]),
    .outData_7(stage_9_per_out[7]),
    .outData_8(stage_9_per_out[8]),
    .outData_9(stage_9_per_out[9]),
    .outData_10(stage_9_per_out[10]),
    .outData_11(stage_9_per_out[11]),
    .outData_12(stage_9_per_out[12]),
    .outData_13(stage_9_per_out[13]),
    .outData_14(stage_9_per_out[14]),
    .outData_15(stage_9_per_out[15]),
    .outData_16(stage_9_per_out[16]),
    .outData_17(stage_9_per_out[17]),
    .outData_18(stage_9_per_out[18]),
    .outData_19(stage_9_per_out[19]),
    .outData_20(stage_9_per_out[20]),
    .outData_21(stage_9_per_out[21]),
    .outData_22(stage_9_per_out[22]),
    .outData_23(stage_9_per_out[23]),
    .outData_24(stage_9_per_out[24]),
    .outData_25(stage_9_per_out[25]),
    .outData_26(stage_9_per_out[26]),
    .outData_27(stage_9_per_out[27]),
    .outData_28(stage_9_per_out[28]),
    .outData_29(stage_9_per_out[29]),
    .outData_30(stage_9_per_out[30]),
    .outData_31(stage_9_per_out[31]),
    .in_start(in_start[9]),
    .out_start(out_start[9]),
    .clk(clk),
    .rst(rst)
  );

  // TODO(Tian): stage 10 32 butterfly units
  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_0 (
    .x_in(stage_9_per_out[0]),
    .y_in(stage_9_per_out[1]),
    .x_out(stage_10_per_in[0]),
    .y_out(stage_10_per_in[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_1 (
    .x_in(stage_9_per_out[2]),
    .y_in(stage_9_per_out[3]),
    .x_out(stage_10_per_in[2]),
    .y_out(stage_10_per_in[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_2 (
    .x_in(stage_9_per_out[4]),
    .y_in(stage_9_per_out[5]),
    .x_out(stage_10_per_in[4]),
    .y_out(stage_10_per_in[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_3 (
    .x_in(stage_9_per_out[6]),
    .y_in(stage_9_per_out[7]),
    .x_out(stage_10_per_in[6]),
    .y_out(stage_10_per_in[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_4 (
    .x_in(stage_9_per_out[8]),
    .y_in(stage_9_per_out[9]),
    .x_out(stage_10_per_in[8]),
    .y_out(stage_10_per_in[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_5 (
    .x_in(stage_9_per_out[10]),
    .y_in(stage_9_per_out[11]),
    .x_out(stage_10_per_in[10]),
    .y_out(stage_10_per_in[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_6 (
    .x_in(stage_9_per_out[12]),
    .y_in(stage_9_per_out[13]),
    .x_out(stage_10_per_in[12]),
    .y_out(stage_10_per_in[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_7 (
    .x_in(stage_9_per_out[14]),
    .y_in(stage_9_per_out[15]),
    .x_out(stage_10_per_in[14]),
    .y_out(stage_10_per_in[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_8 (
    .x_in(stage_9_per_out[16]),
    .y_in(stage_9_per_out[17]),
    .x_out(stage_10_per_in[16]),
    .y_out(stage_10_per_in[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_9 (
    .x_in(stage_9_per_out[18]),
    .y_in(stage_9_per_out[19]),
    .x_out(stage_10_per_in[18]),
    .y_out(stage_10_per_in[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_10 (
    .x_in(stage_9_per_out[20]),
    .y_in(stage_9_per_out[21]),
    .x_out(stage_10_per_in[20]),
    .y_out(stage_10_per_in[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_11 (
    .x_in(stage_9_per_out[22]),
    .y_in(stage_9_per_out[23]),
    .x_out(stage_10_per_in[22]),
    .y_out(stage_10_per_in[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_12 (
    .x_in(stage_9_per_out[24]),
    .y_in(stage_9_per_out[25]),
    .x_out(stage_10_per_in[24]),
    .y_out(stage_10_per_in[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_13 (
    .x_in(stage_9_per_out[26]),
    .y_in(stage_9_per_out[27]),
    .x_out(stage_10_per_in[26]),
    .y_out(stage_10_per_in[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_14 (
    .x_in(stage_9_per_out[28]),
    .y_in(stage_9_per_out[29]),
    .x_out(stage_10_per_in[28]),
    .y_out(stage_10_per_in[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[10]),
    .factors({183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802, 183496802,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570,
              185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570, 185593570}))
  stage_10_butterfly_15 (
    .x_in(stage_9_per_out[30]),
    .y_in(stage_9_per_out[31]),
    .x_out(stage_10_per_in[30]),
    .y_out(stage_10_per_in[31]),
    .clk(clk),
    .rst(rst)
  );


  // TODO(Yang): Update stride
  stage_10_permutation //#(
    //.DATA_WIDTH_PER_INPUT(DATA_WIDTH_PER_INPUT),
    //.INPUT_PER_CYCLE(INPUT_PER_CYCLE))
  stage_10_11_per (
    .inData_0(stage_10_per_in[0]),
    .inData_1(stage_10_per_in[1]),
    .inData_2(stage_10_per_in[2]),
    .inData_3(stage_10_per_in[3]),
    .inData_4(stage_10_per_in[4]),
    .inData_5(stage_10_per_in[5]),
    .inData_6(stage_10_per_in[6]),
    .inData_7(stage_10_per_in[7]),
    .inData_8(stage_10_per_in[8]),
    .inData_9(stage_10_per_in[9]),
    .inData_10(stage_10_per_in[10]),
    .inData_11(stage_10_per_in[11]),
    .inData_12(stage_10_per_in[12]),
    .inData_13(stage_10_per_in[13]),
    .inData_14(stage_10_per_in[14]),
    .inData_15(stage_10_per_in[15]),
    .inData_16(stage_10_per_in[16]),
    .inData_17(stage_10_per_in[17]),
    .inData_18(stage_10_per_in[18]),
    .inData_19(stage_10_per_in[19]),
    .inData_20(stage_10_per_in[20]),
    .inData_21(stage_10_per_in[21]),
    .inData_22(stage_10_per_in[22]),
    .inData_23(stage_10_per_in[23]),
    .inData_24(stage_10_per_in[24]),
    .inData_25(stage_10_per_in[25]),
    .inData_26(stage_10_per_in[26]),
    .inData_27(stage_10_per_in[27]),
    .inData_28(stage_10_per_in[28]),
    .inData_29(stage_10_per_in[29]),
    .inData_30(stage_10_per_in[30]),
    .inData_31(stage_10_per_in[31]),
    .outData_0(stage_10_per_out[0]),
    .outData_1(stage_10_per_out[1]),
    .outData_2(stage_10_per_out[2]),
    .outData_3(stage_10_per_out[3]),
    .outData_4(stage_10_per_out[4]),
    .outData_5(stage_10_per_out[5]),
    .outData_6(stage_10_per_out[6]),
    .outData_7(stage_10_per_out[7]),
    .outData_8(stage_10_per_out[8]),
    .outData_9(stage_10_per_out[9]),
    .outData_10(stage_10_per_out[10]),
    .outData_11(stage_10_per_out[11]),
    .outData_12(stage_10_per_out[12]),
    .outData_13(stage_10_per_out[13]),
    .outData_14(stage_10_per_out[14]),
    .outData_15(stage_10_per_out[15]),
    .outData_16(stage_10_per_out[16]),
    .outData_17(stage_10_per_out[17]),
    .outData_18(stage_10_per_out[18]),
    .outData_19(stage_10_per_out[19]),
    .outData_20(stage_10_per_out[20]),
    .outData_21(stage_10_per_out[21]),
    .outData_22(stage_10_per_out[22]),
    .outData_23(stage_10_per_out[23]),
    .outData_24(stage_10_per_out[24]),
    .outData_25(stage_10_per_out[25]),
    .outData_26(stage_10_per_out[26]),
    .outData_27(stage_10_per_out[27]),
    .outData_28(stage_10_per_out[28]),
    .outData_29(stage_10_per_out[29]),
    .outData_30(stage_10_per_out[30]),
    .outData_31(stage_10_per_out[31]),
    .in_start(in_start[10]),
    .out_start(out_start[10]),
    .clk(clk),
    .rst(rst)
  );

  // TODO(Tian): stage 11 32 butterfly units
  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_0 (
    .x_in(stage_10_per_out[0]),
    .y_in(stage_10_per_out[1]),
    .x_out(outData[0]),
    .y_out(outData[1]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_1 (
    .x_in(stage_10_per_out[2]),
    .y_in(stage_10_per_out[3]),
    .x_out(outData[2]),
    .y_out(outData[3]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_2 (
    .x_in(stage_10_per_out[4]),
    .y_in(stage_10_per_out[5]),
    .x_out(outData[4]),
    .y_out(outData[5]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_3 (
    .x_in(stage_10_per_out[6]),
    .y_in(stage_10_per_out[7]),
    .x_out(outData[6]),
    .y_out(outData[7]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_4 (
    .x_in(stage_10_per_out[8]),
    .y_in(stage_10_per_out[9]),
    .x_out(outData[8]),
    .y_out(outData[9]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_5 (
    .x_in(stage_10_per_out[10]),
    .y_in(stage_10_per_out[11]),
    .x_out(outData[10]),
    .y_out(outData[11]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_6 (
    .x_in(stage_10_per_out[12]),
    .y_in(stage_10_per_out[13]),
    .x_out(outData[12]),
    .y_out(outData[13]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_7 (
    .x_in(stage_10_per_out[14]),
    .y_in(stage_10_per_out[15]),
    .x_out(outData[14]),
    .y_out(outData[15]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_8 (
    .x_in(stage_10_per_out[16]),
    .y_in(stage_10_per_out[17]),
    .x_out(outData[16]),
    .y_out(outData[17]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_9 (
    .x_in(stage_10_per_out[18]),
    .y_in(stage_10_per_out[19]),
    .x_out(outData[18]),
    .y_out(outData[19]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_10 (
    .x_in(stage_10_per_out[20]),
    .y_in(stage_10_per_out[21]),
    .x_out(outData[20]),
    .y_out(outData[21]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_11 (
    .x_in(stage_10_per_out[22]),
    .y_in(stage_10_per_out[23]),
    .x_out(outData[22]),
    .y_out(outData[23]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_12 (
    .x_in(stage_10_per_out[24]),
    .y_in(stage_10_per_out[25]),
    .x_out(outData[24]),
    .y_out(outData[25]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_13 (
    .x_in(stage_10_per_out[26]),
    .y_in(stage_10_per_out[27]),
    .x_out(outData[26]),
    .y_out(outData[27]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_14 (
    .x_in(stage_10_per_out[28]),
    .y_in(stage_10_per_out[29]),
    .x_out(outData[28]),
    .y_out(outData[29]),
    .clk(clk),
    .rst(rst)
  );

  butterfly #(
    .start(START_CYCLE[11]),
    .factors({193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160,
              193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160, 193295160}))
  stage_11_butterfly_15 (
    .x_in(stage_10_per_out[30]),
    .y_in(stage_10_per_out[31]),
    .x_out(outData[30]),
    .y_out(outData[31]),
    .clk(clk),
    .rst(rst)
  );



endmodule
